module aes_128(clk, state, key, out);

    input         clk;
    input  [127:0] state, key;
    output [127:0] out;
				   
    reg [7:0]   p00, p01, p02, p03,
                p10, p11, p12, p13,
                p20, p21, p22, p23,
                p30, p31, p32, p33;
				
    reg [31:0] k0, k1, k2, k3;

    wire [31:0]  s0, s1, s2, s3,
                 z0, z1, z2, z3;

    assign {s0, s1, s2, s3} = state ^ key;
	
    always @ (posedge clk)

    begin
	
    {k0, k1, k2, k3} = key;
	
	// **************************** PART S0 ****************************
	
    // First Portion
    case (s0[7:0])
    8'h00: p00 <= 8'h63;
    8'h01: p00 <= 8'h7c;
    8'h02: p00 <= 8'h77;
    8'h03: p00 <= 8'h7b;
    8'h04: p00 <= 8'hf2;
    8'h05: p00 <= 8'h6b;
    8'h06: p00 <= 8'h6f;
    8'h07: p00 <= 8'hc5;
    8'h08: p00 <= 8'h30;
    8'h09: p00 <= 8'h01;
    8'h0a: p00 <= 8'h67;
    8'h0b: p00 <= 8'h2b;
    8'h0c: p00 <= 8'hfe;
    8'h0d: p00 <= 8'hd7;
    8'h0e: p00 <= 8'hab;
    8'h0f: p00 <= 8'h76;
    8'h10: p00 <= 8'hca;
    8'h11: p00 <= 8'h82;
    8'h12: p00 <= 8'hc9;
    8'h13: p00 <= 8'h7d;
    8'h14: p00 <= 8'hfa;
    8'h15: p00 <= 8'h59;
    8'h16: p00 <= 8'h47;
    8'h17: p00 <= 8'hf0;
    8'h18: p00 <= 8'had;
    8'h19: p00 <= 8'hd4;
    8'h1a: p00 <= 8'ha2;
    8'h1b: p00 <= 8'haf;
    8'h1c: p00 <= 8'h9c;
    8'h1d: p00 <= 8'ha4;
    8'h1e: p00 <= 8'h72;
    8'h1f: p00 <= 8'hc0;
    8'h20: p00 <= 8'hb7;
    8'h21: p00 <= 8'hfd;
    8'h22: p00 <= 8'h93;
    8'h23: p00 <= 8'h26;
    8'h24: p00 <= 8'h36;
    8'h25: p00 <= 8'h3f;
    8'h26: p00 <= 8'hf7;
    8'h27: p00 <= 8'hcc;
    8'h28: p00 <= 8'h34;
    8'h29: p00 <= 8'ha5;
    8'h2a: p00 <= 8'he5;
    8'h2b: p00 <= 8'hf1;
    8'h2c: p00 <= 8'h71;
    8'h2d: p00 <= 8'hd8;
    8'h2e: p00 <= 8'h31;
    8'h2f: p00 <= 8'h15;
    8'h30: p00 <= 8'h04;
    8'h31: p00 <= 8'hc7;
    8'h32: p00 <= 8'h23;
    8'h33: p00 <= 8'hc3;
    8'h34: p00 <= 8'h18;
    8'h35: p00 <= 8'h96;
    8'h36: p00 <= 8'h05;
    8'h37: p00 <= 8'h9a;
    8'h38: p00 <= 8'h07;
    8'h39: p00 <= 8'h12;
    8'h3a: p00 <= 8'h80;
    8'h3b: p00 <= 8'he2;
    8'h3c: p00 <= 8'heb;
    8'h3d: p00 <= 8'h27;
    8'h3e: p00 <= 8'hb2;
    8'h3f: p00 <= 8'h75;
    8'h40: p00 <= 8'h09;
    8'h41: p00 <= 8'h83;
    8'h42: p00 <= 8'h2c;
    8'h43: p00 <= 8'h1a;
    8'h44: p00 <= 8'h1b;
    8'h45: p00 <= 8'h6e;
    8'h46: p00 <= 8'h5a;
    8'h47: p00 <= 8'ha0;
    8'h48: p00 <= 8'h52;
    8'h49: p00 <= 8'h3b;
    8'h4a: p00 <= 8'hd6;
    8'h4b: p00 <= 8'hb3;
    8'h4c: p00 <= 8'h29;
    8'h4d: p00 <= 8'he3;
    8'h4e: p00 <= 8'h2f;
    8'h4f: p00 <= 8'h84;
    8'h50: p00 <= 8'h53;
    8'h51: p00 <= 8'hd1;
    8'h52: p00 <= 8'h00;
    8'h53: p00 <= 8'hed;
    8'h54: p00 <= 8'h20;
    8'h55: p00 <= 8'hfc;
    8'h56: p00 <= 8'hb1;
    8'h57: p00 <= 8'h5b;
    8'h58: p00 <= 8'h6a;
    8'h59: p00 <= 8'hcb;
    8'h5a: p00 <= 8'hbe;
    8'h5b: p00 <= 8'h39;
    8'h5c: p00 <= 8'h4a;
    8'h5d: p00 <= 8'h4c;
    8'h5e: p00 <= 8'h58;
    8'h5f: p00 <= 8'hcf;
    8'h60: p00 <= 8'hd0;
    8'h61: p00 <= 8'hef;
    8'h62: p00 <= 8'haa;
    8'h63: p00 <= 8'hfb;
    8'h64: p00 <= 8'h43;
    8'h65: p00 <= 8'h4d;
    8'h66: p00 <= 8'h33;
    8'h67: p00 <= 8'h85;
    8'h68: p00 <= 8'h45;
    8'h69: p00 <= 8'hf9;
    8'h6a: p00 <= 8'h02;
    8'h6b: p00 <= 8'h7f;
    8'h6c: p00 <= 8'h50;
    8'h6d: p00 <= 8'h3c;
    8'h6e: p00 <= 8'h9f;
    8'h6f: p00 <= 8'ha8;
    8'h70: p00 <= 8'h51;
    8'h71: p00 <= 8'ha3;
    8'h72: p00 <= 8'h40;
    8'h73: p00 <= 8'h8f;
    8'h74: p00 <= 8'h92;
    8'h75: p00 <= 8'h9d;
    8'h76: p00 <= 8'h38;
    8'h77: p00 <= 8'hf5;
    8'h78: p00 <= 8'hbc;
    8'h79: p00 <= 8'hb6;
    8'h7a: p00 <= 8'hda;
    8'h7b: p00 <= 8'h21;
    8'h7c: p00 <= 8'h10;
    8'h7d: p00 <= 8'hff;
    8'h7e: p00 <= 8'hf3;
    8'h7f: p00 <= 8'hd2;
    8'h80: p00 <= 8'hcd;
    8'h81: p00 <= 8'h0c;
    8'h82: p00 <= 8'h13;
    8'h83: p00 <= 8'hec;
    8'h84: p00 <= 8'h5f;
    8'h85: p00 <= 8'h97;
    8'h86: p00 <= 8'h44;
    8'h87: p00 <= 8'h17;
    8'h88: p00 <= 8'hc4;
    8'h89: p00 <= 8'ha7;
    8'h8a: p00 <= 8'h7e;
    8'h8b: p00 <= 8'h3d;
    8'h8c: p00 <= 8'h64;
    8'h8d: p00 <= 8'h5d;
    8'h8e: p00 <= 8'h19;
    8'h8f: p00 <= 8'h73;
    8'h90: p00 <= 8'h60;
    8'h91: p00 <= 8'h81;
    8'h92: p00 <= 8'h4f;
    8'h93: p00 <= 8'hdc;
    8'h94: p00 <= 8'h22;
    8'h95: p00 <= 8'h2a;
    8'h96: p00 <= 8'h90;
    8'h97: p00 <= 8'h88;
    8'h98: p00 <= 8'h46;
    8'h99: p00 <= 8'hee;
    8'h9a: p00 <= 8'hb8;
    8'h9b: p00 <= 8'h14;
    8'h9c: p00 <= 8'hde;
    8'h9d: p00 <= 8'h5e;
    8'h9e: p00 <= 8'h0b;
    8'h9f: p00 <= 8'hdb;
    8'ha0: p00 <= 8'he0;
    8'ha1: p00 <= 8'h32;
    8'ha2: p00 <= 8'h3a;
    8'ha3: p00 <= 8'h0a;
    8'ha4: p00 <= 8'h49;
    8'ha5: p00 <= 8'h06;
    8'ha6: p00 <= 8'h24;
    8'ha7: p00 <= 8'h5c;
    8'ha8: p00 <= 8'hc2;
    8'ha9: p00 <= 8'hd3;
    8'haa: p00 <= 8'hac;
    8'hab: p00 <= 8'h62;
    8'hac: p00 <= 8'h91;
    8'had: p00 <= 8'h95;
    8'hae: p00 <= 8'he4;
    8'haf: p00 <= 8'h79;
    8'hb0: p00 <= 8'he7;
    8'hb1: p00 <= 8'hc8;
    8'hb2: p00 <= 8'h37;
    8'hb3: p00 <= 8'h6d;
    8'hb4: p00 <= 8'h8d;
    8'hb5: p00 <= 8'hd5;
    8'hb6: p00 <= 8'h4e;
    8'hb7: p00 <= 8'ha9;
    8'hb8: p00 <= 8'h6c;
    8'hb9: p00 <= 8'h56;
    8'hba: p00 <= 8'hf4;
    8'hbb: p00 <= 8'hea;
    8'hbc: p00 <= 8'h65;
    8'hbd: p00 <= 8'h7a;
    8'hbe: p00 <= 8'hae;
    8'hbf: p00 <= 8'h08;
    8'hc0: p00 <= 8'hba;
    8'hc1: p00 <= 8'h78;
    8'hc2: p00 <= 8'h25;
    8'hc3: p00 <= 8'h2e;
    8'hc4: p00 <= 8'h1c;
    8'hc5: p00 <= 8'ha6;
    8'hc6: p00 <= 8'hb4;
    8'hc7: p00 <= 8'hc6;
    8'hc8: p00 <= 8'he8;
    8'hc9: p00 <= 8'hdd;
    8'hca: p00 <= 8'h74;
    8'hcb: p00 <= 8'h1f;
    8'hcc: p00 <= 8'h4b;
    8'hcd: p00 <= 8'hbd;
    8'hce: p00 <= 8'h8b;
    8'hcf: p00 <= 8'h8a;
    8'hd0: p00 <= 8'h70;
    8'hd1: p00 <= 8'h3e;
    8'hd2: p00 <= 8'hb5;
    8'hd3: p00 <= 8'h66;
    8'hd4: p00 <= 8'h48;
    8'hd5: p00 <= 8'h03;
    8'hd6: p00 <= 8'hf6;
    8'hd7: p00 <= 8'h0e;
    8'hd8: p00 <= 8'h61;
    8'hd9: p00 <= 8'h35;
    8'hda: p00 <= 8'h57;
    8'hdb: p00 <= 8'hb9;
    8'hdc: p00 <= 8'h86;
    8'hdd: p00 <= 8'hc1;
    8'hde: p00 <= 8'h1d;
    8'hdf: p00 <= 8'h9e;
    8'he0: p00 <= 8'he1;
    8'he1: p00 <= 8'hf8;
    8'he2: p00 <= 8'h98;
    8'he3: p00 <= 8'h11;
    8'he4: p00 <= 8'h69;
    8'he5: p00 <= 8'hd9;
    8'he6: p00 <= 8'h8e;
    8'he7: p00 <= 8'h94;
    8'he8: p00 <= 8'h9b;
    8'he9: p00 <= 8'h1e;
    8'hea: p00 <= 8'h87;
    8'heb: p00 <= 8'he9;
    8'hec: p00 <= 8'hce;
    8'hed: p00 <= 8'h55;
    8'hee: p00 <= 8'h28;
    8'hef: p00 <= 8'hdf;
    8'hf0: p00 <= 8'h8c;
    8'hf1: p00 <= 8'ha1;
    8'hf2: p00 <= 8'h89;
    8'hf3: p00 <= 8'h0d;
    8'hf4: p00 <= 8'hbf;
    8'hf5: p00 <= 8'he6;
    8'hf6: p00 <= 8'h42;
    8'hf7: p00 <= 8'h68;
    8'hf8: p00 <= 8'h41;
    8'hf9: p00 <= 8'h99;
    8'hfa: p00 <= 8'h2d;
    8'hfb: p00 <= 8'h0f;
    8'hfc: p00 <= 8'hb0;
    8'hfd: p00 <= 8'h54;
    8'hfe: p00 <= 8'hbb;
    8'hff: p00 <= 8'h16;
    endcase
	
    // Second Portion
    case (s0[15:8])
    8'h00: p01 <= 8'h63;
    8'h01: p01 <= 8'h7c;
    8'h02: p01 <= 8'h77;
    8'h03: p01 <= 8'h7b;
    8'h04: p01 <= 8'hf2;
    8'h05: p01 <= 8'h6b;
    8'h06: p01 <= 8'h6f;
    8'h07: p01 <= 8'hc5;
    8'h08: p01 <= 8'h30;
    8'h09: p01 <= 8'h01;
    8'h0a: p01 <= 8'h67;
    8'h0b: p01 <= 8'h2b;
    8'h0c: p01 <= 8'hfe;
    8'h0d: p01 <= 8'hd7;
    8'h0e: p01 <= 8'hab;
    8'h0f: p01 <= 8'h76;
    8'h10: p01 <= 8'hca;
    8'h11: p01 <= 8'h82;
    8'h12: p01 <= 8'hc9;
    8'h13: p01 <= 8'h7d;
    8'h14: p01 <= 8'hfa;
    8'h15: p01 <= 8'h59;
    8'h16: p01 <= 8'h47;
    8'h17: p01 <= 8'hf0;
    8'h18: p01 <= 8'had;
    8'h19: p01 <= 8'hd4;
    8'h1a: p01 <= 8'ha2;
    8'h1b: p01 <= 8'haf;
    8'h1c: p01 <= 8'h9c;
    8'h1d: p01 <= 8'ha4;
    8'h1e: p01 <= 8'h72;
    8'h1f: p01 <= 8'hc0;
    8'h20: p01 <= 8'hb7;
    8'h21: p01 <= 8'hfd;
    8'h22: p01 <= 8'h93;
    8'h23: p01 <= 8'h26;
    8'h24: p01 <= 8'h36;
    8'h25: p01 <= 8'h3f;
    8'h26: p01 <= 8'hf7;
    8'h27: p01 <= 8'hcc;
    8'h28: p01 <= 8'h34;
    8'h29: p01 <= 8'ha5;
    8'h2a: p01 <= 8'he5;
    8'h2b: p01 <= 8'hf1;
    8'h2c: p01 <= 8'h71;
    8'h2d: p01 <= 8'hd8;
    8'h2e: p01 <= 8'h31;
    8'h2f: p01 <= 8'h15;
    8'h30: p01 <= 8'h04;
    8'h31: p01 <= 8'hc7;
    8'h32: p01 <= 8'h23;
    8'h33: p01 <= 8'hc3;
    8'h34: p01 <= 8'h18;
    8'h35: p01 <= 8'h96;
    8'h36: p01 <= 8'h05;
    8'h37: p01 <= 8'h9a;
    8'h38: p01 <= 8'h07;
    8'h39: p01 <= 8'h12;
    8'h3a: p01 <= 8'h80;
    8'h3b: p01 <= 8'he2;
    8'h3c: p01 <= 8'heb;
    8'h3d: p01 <= 8'h27;
    8'h3e: p01 <= 8'hb2;
    8'h3f: p01 <= 8'h75;
    8'h40: p01 <= 8'h09;
    8'h41: p01 <= 8'h83;
    8'h42: p01 <= 8'h2c;
    8'h43: p01 <= 8'h1a;
    8'h44: p01 <= 8'h1b;
    8'h45: p01 <= 8'h6e;
    8'h46: p01 <= 8'h5a;
    8'h47: p01 <= 8'ha0;
    8'h48: p01 <= 8'h52;
    8'h49: p01 <= 8'h3b;
    8'h4a: p01 <= 8'hd6;
    8'h4b: p01 <= 8'hb3;
    8'h4c: p01 <= 8'h29;
    8'h4d: p01 <= 8'he3;
    8'h4e: p01 <= 8'h2f;
    8'h4f: p01 <= 8'h84;
    8'h50: p01 <= 8'h53;
    8'h51: p01 <= 8'hd1;
    8'h52: p01 <= 8'h00;
    8'h53: p01 <= 8'hed;
    8'h54: p01 <= 8'h20;
    8'h55: p01 <= 8'hfc;
    8'h56: p01 <= 8'hb1;
    8'h57: p01 <= 8'h5b;
    8'h58: p01 <= 8'h6a;
    8'h59: p01 <= 8'hcb;
    8'h5a: p01 <= 8'hbe;
    8'h5b: p01 <= 8'h39;
    8'h5c: p01 <= 8'h4a;
    8'h5d: p01 <= 8'h4c;
    8'h5e: p01 <= 8'h58;
    8'h5f: p01 <= 8'hcf;
    8'h60: p01 <= 8'hd0;
    8'h61: p01 <= 8'hef;
    8'h62: p01 <= 8'haa;
    8'h63: p01 <= 8'hfb;
    8'h64: p01 <= 8'h43;
    8'h65: p01 <= 8'h4d;
    8'h66: p01 <= 8'h33;
    8'h67: p01 <= 8'h85;
    8'h68: p01 <= 8'h45;
    8'h69: p01 <= 8'hf9;
    8'h6a: p01 <= 8'h02;
    8'h6b: p01 <= 8'h7f;
    8'h6c: p01 <= 8'h50;
    8'h6d: p01 <= 8'h3c;
    8'h6e: p01 <= 8'h9f;
    8'h6f: p01 <= 8'ha8;
    8'h70: p01 <= 8'h51;
    8'h71: p01 <= 8'ha3;
    8'h72: p01 <= 8'h40;
    8'h73: p01 <= 8'h8f;
    8'h74: p01 <= 8'h92;
    8'h75: p01 <= 8'h9d;
    8'h76: p01 <= 8'h38;
    8'h77: p01 <= 8'hf5;
    8'h78: p01 <= 8'hbc;
    8'h79: p01 <= 8'hb6;
    8'h7a: p01 <= 8'hda;
    8'h7b: p01 <= 8'h21;
    8'h7c: p01 <= 8'h10;
    8'h7d: p01 <= 8'hff;
    8'h7e: p01 <= 8'hf3;
    8'h7f: p01 <= 8'hd2;
    8'h80: p01 <= 8'hcd;
    8'h81: p01 <= 8'h0c;
    8'h82: p01 <= 8'h13;
    8'h83: p01 <= 8'hec;
    8'h84: p01 <= 8'h5f;
    8'h85: p01 <= 8'h97;
    8'h86: p01 <= 8'h44;
    8'h87: p01 <= 8'h17;
    8'h88: p01 <= 8'hc4;
    8'h89: p01 <= 8'ha7;
    8'h8a: p01 <= 8'h7e;
    8'h8b: p01 <= 8'h3d;
    8'h8c: p01 <= 8'h64;
    8'h8d: p01 <= 8'h5d;
    8'h8e: p01 <= 8'h19;
    8'h8f: p01 <= 8'h73;
    8'h90: p01 <= 8'h60;
    8'h91: p01 <= 8'h81;
    8'h92: p01 <= 8'h4f;
    8'h93: p01 <= 8'hdc;
    8'h94: p01 <= 8'h22;
    8'h95: p01 <= 8'h2a;
    8'h96: p01 <= 8'h90;
    8'h97: p01 <= 8'h88;
    8'h98: p01 <= 8'h46;
    8'h99: p01 <= 8'hee;
    8'h9a: p01 <= 8'hb8;
    8'h9b: p01 <= 8'h14;
    8'h9c: p01 <= 8'hde;
    8'h9d: p01 <= 8'h5e;
    8'h9e: p01 <= 8'h0b;
    8'h9f: p01 <= 8'hdb;
    8'ha0: p01 <= 8'he0;
    8'ha1: p01 <= 8'h32;
    8'ha2: p01 <= 8'h3a;
    8'ha3: p01 <= 8'h0a;
    8'ha4: p01 <= 8'h49;
    8'ha5: p01 <= 8'h06;
    8'ha6: p01 <= 8'h24;
    8'ha7: p01 <= 8'h5c;
    8'ha8: p01 <= 8'hc2;
    8'ha9: p01 <= 8'hd3;
    8'haa: p01 <= 8'hac;
    8'hab: p01 <= 8'h62;
    8'hac: p01 <= 8'h91;
    8'had: p01 <= 8'h95;
    8'hae: p01 <= 8'he4;
    8'haf: p01 <= 8'h79;
    8'hb0: p01 <= 8'he7;
    8'hb1: p01 <= 8'hc8;
    8'hb2: p01 <= 8'h37;
    8'hb3: p01 <= 8'h6d;
    8'hb4: p01 <= 8'h8d;
    8'hb5: p01 <= 8'hd5;
    8'hb6: p01 <= 8'h4e;
    8'hb7: p01 <= 8'ha9;
    8'hb8: p01 <= 8'h6c;
    8'hb9: p01 <= 8'h56;
    8'hba: p01 <= 8'hf4;
    8'hbb: p01 <= 8'hea;
    8'hbc: p01 <= 8'h65;
    8'hbd: p01 <= 8'h7a;
    8'hbe: p01 <= 8'hae;
    8'hbf: p01 <= 8'h08;
    8'hc0: p01 <= 8'hba;
    8'hc1: p01 <= 8'h78;
    8'hc2: p01 <= 8'h25;
    8'hc3: p01 <= 8'h2e;
    8'hc4: p01 <= 8'h1c;
    8'hc5: p01 <= 8'ha6;
    8'hc6: p01 <= 8'hb4;
    8'hc7: p01 <= 8'hc6;
    8'hc8: p01 <= 8'he8;
    8'hc9: p01 <= 8'hdd;
    8'hca: p01 <= 8'h74;
    8'hcb: p01 <= 8'h1f;
    8'hcc: p01 <= 8'h4b;
    8'hcd: p01 <= 8'hbd;
    8'hce: p01 <= 8'h8b;
    8'hcf: p01 <= 8'h8a;
    8'hd0: p01 <= 8'h70;
    8'hd1: p01 <= 8'h3e;
    8'hd2: p01 <= 8'hb5;
    8'hd3: p01 <= 8'h66;
    8'hd4: p01 <= 8'h48;
    8'hd5: p01 <= 8'h03;
    8'hd6: p01 <= 8'hf6;
    8'hd7: p01 <= 8'h0e;
    8'hd8: p01 <= 8'h61;
    8'hd9: p01 <= 8'h35;
    8'hda: p01 <= 8'h57;
    8'hdb: p01 <= 8'hb9;
    8'hdc: p01 <= 8'h86;
    8'hdd: p01 <= 8'hc1;
    8'hde: p01 <= 8'h1d;
    8'hdf: p01 <= 8'h9e;
    8'he0: p01 <= 8'he1;
    8'he1: p01 <= 8'hf8;
    8'he2: p01 <= 8'h98;
    8'he3: p01 <= 8'h11;
    8'he4: p01 <= 8'h69;
    8'he5: p01 <= 8'hd9;
    8'he6: p01 <= 8'h8e;
    8'he7: p01 <= 8'h94;
    8'he8: p01 <= 8'h9b;
    8'he9: p01 <= 8'h1e;
    8'hea: p01 <= 8'h87;
    8'heb: p01 <= 8'he9;
    8'hec: p01 <= 8'hce;
    8'hed: p01 <= 8'h55;
    8'hee: p01 <= 8'h28;
    8'hef: p01 <= 8'hdf;
    8'hf0: p01 <= 8'h8c;
    8'hf1: p01 <= 8'ha1;
    8'hf2: p01 <= 8'h89;
    8'hf3: p01 <= 8'h0d;
    8'hf4: p01 <= 8'hbf;
    8'hf5: p01 <= 8'he6;
    8'hf6: p01 <= 8'h42;
    8'hf7: p01 <= 8'h68;
    8'hf8: p01 <= 8'h41;
    8'hf9: p01 <= 8'h99;
    8'hfa: p01 <= 8'h2d;
    8'hfb: p01 <= 8'h0f;
    8'hfc: p01 <= 8'hb0;
    8'hfd: p01 <= 8'h54;
    8'hfe: p01 <= 8'hbb;
    8'hff: p01 <= 8'h16;
    endcase
	
    // Third Portion
    case (s0[23:16])
    8'h00: p02 <= 8'h63;
    8'h01: p02 <= 8'h7c;
    8'h02: p02 <= 8'h77;
    8'h03: p02 <= 8'h7b;
    8'h04: p02 <= 8'hf2;
    8'h05: p02 <= 8'h6b;
    8'h06: p02 <= 8'h6f;
    8'h07: p02 <= 8'hc5;
    8'h08: p02 <= 8'h30;
    8'h09: p02 <= 8'h01;
    8'h0a: p02 <= 8'h67;
    8'h0b: p02 <= 8'h2b;
    8'h0c: p02 <= 8'hfe;
    8'h0d: p02 <= 8'hd7;
    8'h0e: p02 <= 8'hab;
    8'h0f: p02 <= 8'h76;
    8'h10: p02 <= 8'hca;
    8'h11: p02 <= 8'h82;
    8'h12: p02 <= 8'hc9;
    8'h13: p02 <= 8'h7d;
    8'h14: p02 <= 8'hfa;
    8'h15: p02 <= 8'h59;
    8'h16: p02 <= 8'h47;
    8'h17: p02 <= 8'hf0;
    8'h18: p02 <= 8'had;
    8'h19: p02 <= 8'hd4;
    8'h1a: p02 <= 8'ha2;
    8'h1b: p02 <= 8'haf;
    8'h1c: p02 <= 8'h9c;
    8'h1d: p02 <= 8'ha4;
    8'h1e: p02 <= 8'h72;
    8'h1f: p02 <= 8'hc0;
    8'h20: p02 <= 8'hb7;
    8'h21: p02 <= 8'hfd;
    8'h22: p02 <= 8'h93;
    8'h23: p02 <= 8'h26;
    8'h24: p02 <= 8'h36;
    8'h25: p02 <= 8'h3f;
    8'h26: p02 <= 8'hf7;
    8'h27: p02 <= 8'hcc;
    8'h28: p02 <= 8'h34;
    8'h29: p02 <= 8'ha5;
    8'h2a: p02 <= 8'he5;
    8'h2b: p02 <= 8'hf1;
    8'h2c: p02 <= 8'h71;
    8'h2d: p02 <= 8'hd8;
    8'h2e: p02 <= 8'h31;
    8'h2f: p02 <= 8'h15;
    8'h30: p02 <= 8'h04;
    8'h31: p02 <= 8'hc7;
    8'h32: p02 <= 8'h23;
    8'h33: p02 <= 8'hc3;
    8'h34: p02 <= 8'h18;
    8'h35: p02 <= 8'h96;
    8'h36: p02 <= 8'h05;
    8'h37: p02 <= 8'h9a;
    8'h38: p02 <= 8'h07;
    8'h39: p02 <= 8'h12;
    8'h3a: p02 <= 8'h80;
    8'h3b: p02 <= 8'he2;
    8'h3c: p02 <= 8'heb;
    8'h3d: p02 <= 8'h27;
    8'h3e: p02 <= 8'hb2;
    8'h3f: p02 <= 8'h75;
    8'h40: p02 <= 8'h09;
    8'h41: p02 <= 8'h83;
    8'h42: p02 <= 8'h2c;
    8'h43: p02 <= 8'h1a;
    8'h44: p02 <= 8'h1b;
    8'h45: p02 <= 8'h6e;
    8'h46: p02 <= 8'h5a;
    8'h47: p02 <= 8'ha0;
    8'h48: p02 <= 8'h52;
    8'h49: p02 <= 8'h3b;
    8'h4a: p02 <= 8'hd6;
    8'h4b: p02 <= 8'hb3;
    8'h4c: p02 <= 8'h29;
    8'h4d: p02 <= 8'he3;
    8'h4e: p02 <= 8'h2f;
    8'h4f: p02 <= 8'h84;
    8'h50: p02 <= 8'h53;
    8'h51: p02 <= 8'hd1;
    8'h52: p02 <= 8'h00;
    8'h53: p02 <= 8'hed;
    8'h54: p02 <= 8'h20;
    8'h55: p02 <= 8'hfc;
    8'h56: p02 <= 8'hb1;
    8'h57: p02 <= 8'h5b;
    8'h58: p02 <= 8'h6a;
    8'h59: p02 <= 8'hcb;
    8'h5a: p02 <= 8'hbe;
    8'h5b: p02 <= 8'h39;
    8'h5c: p02 <= 8'h4a;
    8'h5d: p02 <= 8'h4c;
    8'h5e: p02 <= 8'h58;
    8'h5f: p02 <= 8'hcf;
    8'h60: p02 <= 8'hd0;
    8'h61: p02 <= 8'hef;
    8'h62: p02 <= 8'haa;
    8'h63: p02 <= 8'hfb;
    8'h64: p02 <= 8'h43;
    8'h65: p02 <= 8'h4d;
    8'h66: p02 <= 8'h33;
    8'h67: p02 <= 8'h85;
    8'h68: p02 <= 8'h45;
    8'h69: p02 <= 8'hf9;
    8'h6a: p02 <= 8'h02;
    8'h6b: p02 <= 8'h7f;
    8'h6c: p02 <= 8'h50;
    8'h6d: p02 <= 8'h3c;
    8'h6e: p02 <= 8'h9f;
    8'h6f: p02 <= 8'ha8;
    8'h70: p02 <= 8'h51;
    8'h71: p02 <= 8'ha3;
    8'h72: p02 <= 8'h40;
    8'h73: p02 <= 8'h8f;
    8'h74: p02 <= 8'h92;
    8'h75: p02 <= 8'h9d;
    8'h76: p02 <= 8'h38;
    8'h77: p02 <= 8'hf5;
    8'h78: p02 <= 8'hbc;
    8'h79: p02 <= 8'hb6;
    8'h7a: p02 <= 8'hda;
    8'h7b: p02 <= 8'h21;
    8'h7c: p02 <= 8'h10;
    8'h7d: p02 <= 8'hff;
    8'h7e: p02 <= 8'hf3;
    8'h7f: p02 <= 8'hd2;
    8'h80: p02 <= 8'hcd;
    8'h81: p02 <= 8'h0c;
    8'h82: p02 <= 8'h13;
    8'h83: p02 <= 8'hec;
    8'h84: p02 <= 8'h5f;
    8'h85: p02 <= 8'h97;
    8'h86: p02 <= 8'h44;
    8'h87: p02 <= 8'h17;
    8'h88: p02 <= 8'hc4;
    8'h89: p02 <= 8'ha7;
    8'h8a: p02 <= 8'h7e;
    8'h8b: p02 <= 8'h3d;
    8'h8c: p02 <= 8'h64;
    8'h8d: p02 <= 8'h5d;
    8'h8e: p02 <= 8'h19;
    8'h8f: p02 <= 8'h73;
    8'h90: p02 <= 8'h60;
    8'h91: p02 <= 8'h81;
    8'h92: p02 <= 8'h4f;
    8'h93: p02 <= 8'hdc;
    8'h94: p02 <= 8'h22;
    8'h95: p02 <= 8'h2a;
    8'h96: p02 <= 8'h90;
    8'h97: p02 <= 8'h88;
    8'h98: p02 <= 8'h46;
    8'h99: p02 <= 8'hee;
    8'h9a: p02 <= 8'hb8;
    8'h9b: p02 <= 8'h14;
    8'h9c: p02 <= 8'hde;
    8'h9d: p02 <= 8'h5e;
    8'h9e: p02 <= 8'h0b;
    8'h9f: p02 <= 8'hdb;
    8'ha0: p02 <= 8'he0;
    8'ha1: p02 <= 8'h32;
    8'ha2: p02 <= 8'h3a;
    8'ha3: p02 <= 8'h0a;
    8'ha4: p02 <= 8'h49;
    8'ha5: p02 <= 8'h06;
    8'ha6: p02 <= 8'h24;
    8'ha7: p02 <= 8'h5c;
    8'ha8: p02 <= 8'hc2;
    8'ha9: p02 <= 8'hd3;
    8'haa: p02 <= 8'hac;
    8'hab: p02 <= 8'h62;
    8'hac: p02 <= 8'h91;
    8'had: p02 <= 8'h95;
    8'hae: p02 <= 8'he4;
    8'haf: p02 <= 8'h79;
    8'hb0: p02 <= 8'he7;
    8'hb1: p02 <= 8'hc8;
    8'hb2: p02 <= 8'h37;
    8'hb3: p02 <= 8'h6d;
    8'hb4: p02 <= 8'h8d;
    8'hb5: p02 <= 8'hd5;
    8'hb6: p02 <= 8'h4e;
    8'hb7: p02 <= 8'ha9;
    8'hb8: p02 <= 8'h6c;
    8'hb9: p02 <= 8'h56;
    8'hba: p02 <= 8'hf4;
    8'hbb: p02 <= 8'hea;
    8'hbc: p02 <= 8'h65;
    8'hbd: p02 <= 8'h7a;
    8'hbe: p02 <= 8'hae;
    8'hbf: p02 <= 8'h08;
    8'hc0: p02 <= 8'hba;
    8'hc1: p02 <= 8'h78;
    8'hc2: p02 <= 8'h25;
    8'hc3: p02 <= 8'h2e;
    8'hc4: p02 <= 8'h1c;
    8'hc5: p02 <= 8'ha6;
    8'hc6: p02 <= 8'hb4;
    8'hc7: p02 <= 8'hc6;
    8'hc8: p02 <= 8'he8;
    8'hc9: p02 <= 8'hdd;
    8'hca: p02 <= 8'h74;
    8'hcb: p02 <= 8'h1f;
    8'hcc: p02 <= 8'h4b;
    8'hcd: p02 <= 8'hbd;
    8'hce: p02 <= 8'h8b;
    8'hcf: p02 <= 8'h8a;
    8'hd0: p02 <= 8'h70;
    8'hd1: p02 <= 8'h3e;
    8'hd2: p02 <= 8'hb5;
    8'hd3: p02 <= 8'h66;
    8'hd4: p02 <= 8'h48;
    8'hd5: p02 <= 8'h03;
    8'hd6: p02 <= 8'hf6;
    8'hd7: p02 <= 8'h0e;
    8'hd8: p02 <= 8'h61;
    8'hd9: p02 <= 8'h35;
    8'hda: p02 <= 8'h57;
    8'hdb: p02 <= 8'hb9;
    8'hdc: p02 <= 8'h86;
    8'hdd: p02 <= 8'hc1;
    8'hde: p02 <= 8'h1d;
    8'hdf: p02 <= 8'h9e;
    8'he0: p02 <= 8'he1;
    8'he1: p02 <= 8'hf8;
    8'he2: p02 <= 8'h98;
    8'he3: p02 <= 8'h11;
    8'he4: p02 <= 8'h69;
    8'he5: p02 <= 8'hd9;
    8'he6: p02 <= 8'h8e;
    8'he7: p02 <= 8'h94;
    8'he8: p02 <= 8'h9b;
    8'he9: p02 <= 8'h1e;
    8'hea: p02 <= 8'h87;
    8'heb: p02 <= 8'he9;
    8'hec: p02 <= 8'hce;
    8'hed: p02 <= 8'h55;
    8'hee: p02 <= 8'h28;
    8'hef: p02 <= 8'hdf;
    8'hf0: p02 <= 8'h8c;
    8'hf1: p02 <= 8'ha1;
    8'hf2: p02 <= 8'h89;
    8'hf3: p02 <= 8'h0d;
    8'hf4: p02 <= 8'hbf;
    8'hf5: p02 <= 8'he6;
    8'hf6: p02 <= 8'h42;
    8'hf7: p02 <= 8'h68;
    8'hf8: p02 <= 8'h41;
    8'hf9: p02 <= 8'h99;
    8'hfa: p02 <= 8'h2d;
    8'hfb: p02 <= 8'h0f;
    8'hfc: p02 <= 8'hb0;
    8'hfd: p02 <= 8'h54;
    8'hfe: p02 <= 8'hbb;
    8'hff: p02 <= 8'h16;
    endcase
	
    // Fourth Portion
    case (s0[31:24])
    8'h00: p03 <= 8'h63;
    8'h01: p03 <= 8'h7c;
    8'h02: p03 <= 8'h77;
    8'h03: p03 <= 8'h7b;
    8'h04: p03 <= 8'hf2;
    8'h05: p03 <= 8'h6b;
    8'h06: p03 <= 8'h6f;
    8'h07: p03 <= 8'hc5;
    8'h08: p03 <= 8'h30;
    8'h09: p03 <= 8'h01;
    8'h0a: p03 <= 8'h67;
    8'h0b: p03 <= 8'h2b;
    8'h0c: p03 <= 8'hfe;
    8'h0d: p03 <= 8'hd7;
    8'h0e: p03 <= 8'hab;
    8'h0f: p03 <= 8'h76;
    8'h10: p03 <= 8'hca;
    8'h11: p03 <= 8'h82;
    8'h12: p03 <= 8'hc9;
    8'h13: p03 <= 8'h7d;
    8'h14: p03 <= 8'hfa;
    8'h15: p03 <= 8'h59;
    8'h16: p03 <= 8'h47;
    8'h17: p03 <= 8'hf0;
    8'h18: p03 <= 8'had;
    8'h19: p03 <= 8'hd4;
    8'h1a: p03 <= 8'ha2;
    8'h1b: p03 <= 8'haf;
    8'h1c: p03 <= 8'h9c;
    8'h1d: p03 <= 8'ha4;
    8'h1e: p03 <= 8'h72;
    8'h1f: p03 <= 8'hc0;
    8'h20: p03 <= 8'hb7;
    8'h21: p03 <= 8'hfd;
    8'h22: p03 <= 8'h93;
    8'h23: p03 <= 8'h26;
    8'h24: p03 <= 8'h36;
    8'h25: p03 <= 8'h3f;
    8'h26: p03 <= 8'hf7;
    8'h27: p03 <= 8'hcc;
    8'h28: p03 <= 8'h34;
    8'h29: p03 <= 8'ha5;
    8'h2a: p03 <= 8'he5;
    8'h2b: p03 <= 8'hf1;
    8'h2c: p03 <= 8'h71;
    8'h2d: p03 <= 8'hd8;
    8'h2e: p03 <= 8'h31;
    8'h2f: p03 <= 8'h15;
    8'h30: p03 <= 8'h04;
    8'h31: p03 <= 8'hc7;
    8'h32: p03 <= 8'h23;
    8'h33: p03 <= 8'hc3;
    8'h34: p03 <= 8'h18;
    8'h35: p03 <= 8'h96;
    8'h36: p03 <= 8'h05;
    8'h37: p03 <= 8'h9a;
    8'h38: p03 <= 8'h07;
    8'h39: p03 <= 8'h12;
    8'h3a: p03 <= 8'h80;
    8'h3b: p03 <= 8'he2;
    8'h3c: p03 <= 8'heb;
    8'h3d: p03 <= 8'h27;
    8'h3e: p03 <= 8'hb2;
    8'h3f: p03 <= 8'h75;
    8'h40: p03 <= 8'h09;
    8'h41: p03 <= 8'h83;
    8'h42: p03 <= 8'h2c;
    8'h43: p03 <= 8'h1a;
    8'h44: p03 <= 8'h1b;
    8'h45: p03 <= 8'h6e;
    8'h46: p03 <= 8'h5a;
    8'h47: p03 <= 8'ha0;
    8'h48: p03 <= 8'h52;
    8'h49: p03 <= 8'h3b;
    8'h4a: p03 <= 8'hd6;
    8'h4b: p03 <= 8'hb3;
    8'h4c: p03 <= 8'h29;
    8'h4d: p03 <= 8'he3;
    8'h4e: p03 <= 8'h2f;
    8'h4f: p03 <= 8'h84;
    8'h50: p03 <= 8'h53;
    8'h51: p03 <= 8'hd1;
    8'h52: p03 <= 8'h00;
    8'h53: p03 <= 8'hed;
    8'h54: p03 <= 8'h20;
    8'h55: p03 <= 8'hfc;
    8'h56: p03 <= 8'hb1;
    8'h57: p03 <= 8'h5b;
    8'h58: p03 <= 8'h6a;
    8'h59: p03 <= 8'hcb;
    8'h5a: p03 <= 8'hbe;
    8'h5b: p03 <= 8'h39;
    8'h5c: p03 <= 8'h4a;
    8'h5d: p03 <= 8'h4c;
    8'h5e: p03 <= 8'h58;
    8'h5f: p03 <= 8'hcf;
    8'h60: p03 <= 8'hd0;
    8'h61: p03 <= 8'hef;
    8'h62: p03 <= 8'haa;
    8'h63: p03 <= 8'hfb;
    8'h64: p03 <= 8'h43;
    8'h65: p03 <= 8'h4d;
    8'h66: p03 <= 8'h33;
    8'h67: p03 <= 8'h85;
    8'h68: p03 <= 8'h45;
    8'h69: p03 <= 8'hf9;
    8'h6a: p03 <= 8'h02;
    8'h6b: p03 <= 8'h7f;
    8'h6c: p03 <= 8'h50;
    8'h6d: p03 <= 8'h3c;
    8'h6e: p03 <= 8'h9f;
    8'h6f: p03 <= 8'ha8;
    8'h70: p03 <= 8'h51;
    8'h71: p03 <= 8'ha3;
    8'h72: p03 <= 8'h40;
    8'h73: p03 <= 8'h8f;
    8'h74: p03 <= 8'h92;
    8'h75: p03 <= 8'h9d;
    8'h76: p03 <= 8'h38;
    8'h77: p03 <= 8'hf5;
    8'h78: p03 <= 8'hbc;
    8'h79: p03 <= 8'hb6;
    8'h7a: p03 <= 8'hda;
    8'h7b: p03 <= 8'h21;
    8'h7c: p03 <= 8'h10;
    8'h7d: p03 <= 8'hff;
    8'h7e: p03 <= 8'hf3;
    8'h7f: p03 <= 8'hd2;
    8'h80: p03 <= 8'hcd;
    8'h81: p03 <= 8'h0c;
    8'h82: p03 <= 8'h13;
    8'h83: p03 <= 8'hec;
    8'h84: p03 <= 8'h5f;
    8'h85: p03 <= 8'h97;
    8'h86: p03 <= 8'h44;
    8'h87: p03 <= 8'h17;
    8'h88: p03 <= 8'hc4;
    8'h89: p03 <= 8'ha7;
    8'h8a: p03 <= 8'h7e;
    8'h8b: p03 <= 8'h3d;
    8'h8c: p03 <= 8'h64;
    8'h8d: p03 <= 8'h5d;
    8'h8e: p03 <= 8'h19;
    8'h8f: p03 <= 8'h73;
    8'h90: p03 <= 8'h60;
    8'h91: p03 <= 8'h81;
    8'h92: p03 <= 8'h4f;
    8'h93: p03 <= 8'hdc;
    8'h94: p03 <= 8'h22;
    8'h95: p03 <= 8'h2a;
    8'h96: p03 <= 8'h90;
    8'h97: p03 <= 8'h88;
    8'h98: p03 <= 8'h46;
    8'h99: p03 <= 8'hee;
    8'h9a: p03 <= 8'hb8;
    8'h9b: p03 <= 8'h14;
    8'h9c: p03 <= 8'hde;
    8'h9d: p03 <= 8'h5e;
    8'h9e: p03 <= 8'h0b;
    8'h9f: p03 <= 8'hdb;
    8'ha0: p03 <= 8'he0;
    8'ha1: p03 <= 8'h32;
    8'ha2: p03 <= 8'h3a;
    8'ha3: p03 <= 8'h0a;
    8'ha4: p03 <= 8'h49;
    8'ha5: p03 <= 8'h06;
    8'ha6: p03 <= 8'h24;
    8'ha7: p03 <= 8'h5c;
    8'ha8: p03 <= 8'hc2;
    8'ha9: p03 <= 8'hd3;
    8'haa: p03 <= 8'hac;
    8'hab: p03 <= 8'h62;
    8'hac: p03 <= 8'h91;
    8'had: p03 <= 8'h95;
    8'hae: p03 <= 8'he4;
    8'haf: p03 <= 8'h79;
    8'hb0: p03 <= 8'he7;
    8'hb1: p03 <= 8'hc8;
    8'hb2: p03 <= 8'h37;
    8'hb3: p03 <= 8'h6d;
    8'hb4: p03 <= 8'h8d;
    8'hb5: p03 <= 8'hd5;
    8'hb6: p03 <= 8'h4e;
    8'hb7: p03 <= 8'ha9;
    8'hb8: p03 <= 8'h6c;
    8'hb9: p03 <= 8'h56;
    8'hba: p03 <= 8'hf4;
    8'hbb: p03 <= 8'hea;
    8'hbc: p03 <= 8'h65;
    8'hbd: p03 <= 8'h7a;
    8'hbe: p03 <= 8'hae;
    8'hbf: p03 <= 8'h08;
    8'hc0: p03 <= 8'hba;
    8'hc1: p03 <= 8'h78;
    8'hc2: p03 <= 8'h25;
    8'hc3: p03 <= 8'h2e;
    8'hc4: p03 <= 8'h1c;
    8'hc5: p03 <= 8'ha6;
    8'hc6: p03 <= 8'hb4;
    8'hc7: p03 <= 8'hc6;
    8'hc8: p03 <= 8'he8;
    8'hc9: p03 <= 8'hdd;
    8'hca: p03 <= 8'h74;
    8'hcb: p03 <= 8'h1f;
    8'hcc: p03 <= 8'h4b;
    8'hcd: p03 <= 8'hbd;
    8'hce: p03 <= 8'h8b;
    8'hcf: p03 <= 8'h8a;
    8'hd0: p03 <= 8'h70;
    8'hd1: p03 <= 8'h3e;
    8'hd2: p03 <= 8'hb5;
    8'hd3: p03 <= 8'h66;
    8'hd4: p03 <= 8'h48;
    8'hd5: p03 <= 8'h03;
    8'hd6: p03 <= 8'hf6;
    8'hd7: p03 <= 8'h0e;
    8'hd8: p03 <= 8'h61;
    8'hd9: p03 <= 8'h35;
    8'hda: p03 <= 8'h57;
    8'hdb: p03 <= 8'hb9;
    8'hdc: p03 <= 8'h86;
    8'hdd: p03 <= 8'hc1;
    8'hde: p03 <= 8'h1d;
    8'hdf: p03 <= 8'h9e;
    8'he0: p03 <= 8'he1;
    8'he1: p03 <= 8'hf8;
    8'he2: p03 <= 8'h98;
    8'he3: p03 <= 8'h11;
    8'he4: p03 <= 8'h69;
    8'he5: p03 <= 8'hd9;
    8'he6: p03 <= 8'h8e;
    8'he7: p03 <= 8'h94;
    8'he8: p03 <= 8'h9b;
    8'he9: p03 <= 8'h1e;
    8'hea: p03 <= 8'h87;
    8'heb: p03 <= 8'he9;
    8'hec: p03 <= 8'hce;
    8'hed: p03 <= 8'h55;
    8'hee: p03 <= 8'h28;
    8'hef: p03 <= 8'hdf;
    8'hf0: p03 <= 8'h8c;
    8'hf1: p03 <= 8'ha1;
    8'hf2: p03 <= 8'h89;
    8'hf3: p03 <= 8'h0d;
    8'hf4: p03 <= 8'hbf;
    8'hf5: p03 <= 8'he6;
    8'hf6: p03 <= 8'h42;
    8'hf7: p03 <= 8'h68;
    8'hf8: p03 <= 8'h41;
    8'hf9: p03 <= 8'h99;
    8'hfa: p03 <= 8'h2d;
    8'hfb: p03 <= 8'h0f;
    8'hfc: p03 <= 8'hb0;
    8'hfd: p03 <= 8'h54;
    8'hfe: p03 <= 8'hbb;
    8'hff: p03 <= 8'h16;
    endcase
	
	// **************************** PART S1 ****************************
	
    // First Portion
    case (s1[7:0])
    8'h00: p10 <= 8'h63;
    8'h01: p10 <= 8'h7c;
    8'h02: p10 <= 8'h77;
    8'h03: p10 <= 8'h7b;
    8'h04: p10 <= 8'hf2;
    8'h05: p10 <= 8'h6b;
    8'h06: p10 <= 8'h6f;
    8'h07: p10 <= 8'hc5;
    8'h08: p10 <= 8'h30;
    8'h09: p10 <= 8'h01;
    8'h0a: p10 <= 8'h67;
    8'h0b: p10 <= 8'h2b;
    8'h0c: p10 <= 8'hfe;
    8'h0d: p10 <= 8'hd7;
    8'h0e: p10 <= 8'hab;
    8'h0f: p10 <= 8'h76;
    8'h10: p10 <= 8'hca;
    8'h11: p10 <= 8'h82;
    8'h12: p10 <= 8'hc9;
    8'h13: p10 <= 8'h7d;
    8'h14: p10 <= 8'hfa;
    8'h15: p10 <= 8'h59;
    8'h16: p10 <= 8'h47;
    8'h17: p10 <= 8'hf0;
    8'h18: p10 <= 8'had;
    8'h19: p10 <= 8'hd4;
    8'h1a: p10 <= 8'ha2;
    8'h1b: p10 <= 8'haf;
    8'h1c: p10 <= 8'h9c;
    8'h1d: p10 <= 8'ha4;
    8'h1e: p10 <= 8'h72;
    8'h1f: p10 <= 8'hc0;
    8'h20: p10 <= 8'hb7;
    8'h21: p10 <= 8'hfd;
    8'h22: p10 <= 8'h93;
    8'h23: p10 <= 8'h26;
    8'h24: p10 <= 8'h36;
    8'h25: p10 <= 8'h3f;
    8'h26: p10 <= 8'hf7;
    8'h27: p10 <= 8'hcc;
    8'h28: p10 <= 8'h34;
    8'h29: p10 <= 8'ha5;
    8'h2a: p10 <= 8'he5;
    8'h2b: p10 <= 8'hf1;
    8'h2c: p10 <= 8'h71;
    8'h2d: p10 <= 8'hd8;
    8'h2e: p10 <= 8'h31;
    8'h2f: p10 <= 8'h15;
    8'h30: p10 <= 8'h04;
    8'h31: p10 <= 8'hc7;
    8'h32: p10 <= 8'h23;
    8'h33: p10 <= 8'hc3;
    8'h34: p10 <= 8'h18;
    8'h35: p10 <= 8'h96;
    8'h36: p10 <= 8'h05;
    8'h37: p10 <= 8'h9a;
    8'h38: p10 <= 8'h07;
    8'h39: p10 <= 8'h12;
    8'h3a: p10 <= 8'h80;
    8'h3b: p10 <= 8'he2;
    8'h3c: p10 <= 8'heb;
    8'h3d: p10 <= 8'h27;
    8'h3e: p10 <= 8'hb2;
    8'h3f: p10 <= 8'h75;
    8'h40: p10 <= 8'h09;
    8'h41: p10 <= 8'h83;
    8'h42: p10 <= 8'h2c;
    8'h43: p10 <= 8'h1a;
    8'h44: p10 <= 8'h1b;
    8'h45: p10 <= 8'h6e;
    8'h46: p10 <= 8'h5a;
    8'h47: p10 <= 8'ha0;
    8'h48: p10 <= 8'h52;
    8'h49: p10 <= 8'h3b;
    8'h4a: p10 <= 8'hd6;
    8'h4b: p10 <= 8'hb3;
    8'h4c: p10 <= 8'h29;
    8'h4d: p10 <= 8'he3;
    8'h4e: p10 <= 8'h2f;
    8'h4f: p10 <= 8'h84;
    8'h50: p10 <= 8'h53;
    8'h51: p10 <= 8'hd1;
    8'h52: p10 <= 8'h00;
    8'h53: p10 <= 8'hed;
    8'h54: p10 <= 8'h20;
    8'h55: p10 <= 8'hfc;
    8'h56: p10 <= 8'hb1;
    8'h57: p10 <= 8'h5b;
    8'h58: p10 <= 8'h6a;
    8'h59: p10 <= 8'hcb;
    8'h5a: p10 <= 8'hbe;
    8'h5b: p10 <= 8'h39;
    8'h5c: p10 <= 8'h4a;
    8'h5d: p10 <= 8'h4c;
    8'h5e: p10 <= 8'h58;
    8'h5f: p10 <= 8'hcf;
    8'h60: p10 <= 8'hd0;
    8'h61: p10 <= 8'hef;
    8'h62: p10 <= 8'haa;
    8'h63: p10 <= 8'hfb;
    8'h64: p10 <= 8'h43;
    8'h65: p10 <= 8'h4d;
    8'h66: p10 <= 8'h33;
    8'h67: p10 <= 8'h85;
    8'h68: p10 <= 8'h45;
    8'h69: p10 <= 8'hf9;
    8'h6a: p10 <= 8'h02;
    8'h6b: p10 <= 8'h7f;
    8'h6c: p10 <= 8'h50;
    8'h6d: p10 <= 8'h3c;
    8'h6e: p10 <= 8'h9f;
    8'h6f: p10 <= 8'ha8;
    8'h70: p10 <= 8'h51;
    8'h71: p10 <= 8'ha3;
    8'h72: p10 <= 8'h40;
    8'h73: p10 <= 8'h8f;
    8'h74: p10 <= 8'h92;
    8'h75: p10 <= 8'h9d;
    8'h76: p10 <= 8'h38;
    8'h77: p10 <= 8'hf5;
    8'h78: p10 <= 8'hbc;
    8'h79: p10 <= 8'hb6;
    8'h7a: p10 <= 8'hda;
    8'h7b: p10 <= 8'h21;
    8'h7c: p10 <= 8'h10;
    8'h7d: p10 <= 8'hff;
    8'h7e: p10 <= 8'hf3;
    8'h7f: p10 <= 8'hd2;
    8'h80: p10 <= 8'hcd;
    8'h81: p10 <= 8'h0c;
    8'h82: p10 <= 8'h13;
    8'h83: p10 <= 8'hec;
    8'h84: p10 <= 8'h5f;
    8'h85: p10 <= 8'h97;
    8'h86: p10 <= 8'h44;
    8'h87: p10 <= 8'h17;
    8'h88: p10 <= 8'hc4;
    8'h89: p10 <= 8'ha7;
    8'h8a: p10 <= 8'h7e;
    8'h8b: p10 <= 8'h3d;
    8'h8c: p10 <= 8'h64;
    8'h8d: p10 <= 8'h5d;
    8'h8e: p10 <= 8'h19;
    8'h8f: p10 <= 8'h73;
    8'h90: p10 <= 8'h60;
    8'h91: p10 <= 8'h81;
    8'h92: p10 <= 8'h4f;
    8'h93: p10 <= 8'hdc;
    8'h94: p10 <= 8'h22;
    8'h95: p10 <= 8'h2a;
    8'h96: p10 <= 8'h90;
    8'h97: p10 <= 8'h88;
    8'h98: p10 <= 8'h46;
    8'h99: p10 <= 8'hee;
    8'h9a: p10 <= 8'hb8;
    8'h9b: p10 <= 8'h14;
    8'h9c: p10 <= 8'hde;
    8'h9d: p10 <= 8'h5e;
    8'h9e: p10 <= 8'h0b;
    8'h9f: p10 <= 8'hdb;
    8'ha0: p10 <= 8'he0;
    8'ha1: p10 <= 8'h32;
    8'ha2: p10 <= 8'h3a;
    8'ha3: p10 <= 8'h0a;
    8'ha4: p10 <= 8'h49;
    8'ha5: p10 <= 8'h06;
    8'ha6: p10 <= 8'h24;
    8'ha7: p10 <= 8'h5c;
    8'ha8: p10 <= 8'hc2;
    8'ha9: p10 <= 8'hd3;
    8'haa: p10 <= 8'hac;
    8'hab: p10 <= 8'h62;
    8'hac: p10 <= 8'h91;
    8'had: p10 <= 8'h95;
    8'hae: p10 <= 8'he4;
    8'haf: p10 <= 8'h79;
    8'hb0: p10 <= 8'he7;
    8'hb1: p10 <= 8'hc8;
    8'hb2: p10 <= 8'h37;
    8'hb3: p10 <= 8'h6d;
    8'hb4: p10 <= 8'h8d;
    8'hb5: p10 <= 8'hd5;
    8'hb6: p10 <= 8'h4e;
    8'hb7: p10 <= 8'ha9;
    8'hb8: p10 <= 8'h6c;
    8'hb9: p10 <= 8'h56;
    8'hba: p10 <= 8'hf4;
    8'hbb: p10 <= 8'hea;
    8'hbc: p10 <= 8'h65;
    8'hbd: p10 <= 8'h7a;
    8'hbe: p10 <= 8'hae;
    8'hbf: p10 <= 8'h08;
    8'hc0: p10 <= 8'hba;
    8'hc1: p10 <= 8'h78;
    8'hc2: p10 <= 8'h25;
    8'hc3: p10 <= 8'h2e;
    8'hc4: p10 <= 8'h1c;
    8'hc5: p10 <= 8'ha6;
    8'hc6: p10 <= 8'hb4;
    8'hc7: p10 <= 8'hc6;
    8'hc8: p10 <= 8'he8;
    8'hc9: p10 <= 8'hdd;
    8'hca: p10 <= 8'h74;
    8'hcb: p10 <= 8'h1f;
    8'hcc: p10 <= 8'h4b;
    8'hcd: p10 <= 8'hbd;
    8'hce: p10 <= 8'h8b;
    8'hcf: p10 <= 8'h8a;
    8'hd0: p10 <= 8'h70;
    8'hd1: p10 <= 8'h3e;
    8'hd2: p10 <= 8'hb5;
    8'hd3: p10 <= 8'h66;
    8'hd4: p10 <= 8'h48;
    8'hd5: p10 <= 8'h03;
    8'hd6: p10 <= 8'hf6;
    8'hd7: p10 <= 8'h0e;
    8'hd8: p10 <= 8'h61;
    8'hd9: p10 <= 8'h35;
    8'hda: p10 <= 8'h57;
    8'hdb: p10 <= 8'hb9;
    8'hdc: p10 <= 8'h86;
    8'hdd: p10 <= 8'hc1;
    8'hde: p10 <= 8'h1d;
    8'hdf: p10 <= 8'h9e;
    8'he0: p10 <= 8'he1;
    8'he1: p10 <= 8'hf8;
    8'he2: p10 <= 8'h98;
    8'he3: p10 <= 8'h11;
    8'he4: p10 <= 8'h69;
    8'he5: p10 <= 8'hd9;
    8'he6: p10 <= 8'h8e;
    8'he7: p10 <= 8'h94;
    8'he8: p10 <= 8'h9b;
    8'he9: p10 <= 8'h1e;
    8'hea: p10 <= 8'h87;
    8'heb: p10 <= 8'he9;
    8'hec: p10 <= 8'hce;
    8'hed: p10 <= 8'h55;
    8'hee: p10 <= 8'h28;
    8'hef: p10 <= 8'hdf;
    8'hf0: p10 <= 8'h8c;
    8'hf1: p10 <= 8'ha1;
    8'hf2: p10 <= 8'h89;
    8'hf3: p10 <= 8'h0d;
    8'hf4: p10 <= 8'hbf;
    8'hf5: p10 <= 8'he6;
    8'hf6: p10 <= 8'h42;
    8'hf7: p10 <= 8'h68;
    8'hf8: p10 <= 8'h41;
    8'hf9: p10 <= 8'h99;
    8'hfa: p10 <= 8'h2d;
    8'hfb: p10 <= 8'h0f;
    8'hfc: p10 <= 8'hb0;
    8'hfd: p10 <= 8'h54;
    8'hfe: p10 <= 8'hbb;
    8'hff: p10 <= 8'h16;
    endcase
	
    // Second Portion
    case (s1[15:8])
    8'h00: p11 <= 8'h63;
    8'h01: p11 <= 8'h7c;
    8'h02: p11 <= 8'h77;
    8'h03: p11 <= 8'h7b;
    8'h04: p11 <= 8'hf2;
    8'h05: p11 <= 8'h6b;
    8'h06: p11 <= 8'h6f;
    8'h07: p11 <= 8'hc5;
    8'h08: p11 <= 8'h30;
    8'h09: p11 <= 8'h01;
    8'h0a: p11 <= 8'h67;
    8'h0b: p11 <= 8'h2b;
    8'h0c: p11 <= 8'hfe;
    8'h0d: p11 <= 8'hd7;
    8'h0e: p11 <= 8'hab;
    8'h0f: p11 <= 8'h76;
    8'h10: p11 <= 8'hca;
    8'h11: p11 <= 8'h82;
    8'h12: p11 <= 8'hc9;
    8'h13: p11 <= 8'h7d;
    8'h14: p11 <= 8'hfa;
    8'h15: p11 <= 8'h59;
    8'h16: p11 <= 8'h47;
    8'h17: p11 <= 8'hf0;
    8'h18: p11 <= 8'had;
    8'h19: p11 <= 8'hd4;
    8'h1a: p11 <= 8'ha2;
    8'h1b: p11 <= 8'haf;
    8'h1c: p11 <= 8'h9c;
    8'h1d: p11 <= 8'ha4;
    8'h1e: p11 <= 8'h72;
    8'h1f: p11 <= 8'hc0;
    8'h20: p11 <= 8'hb7;
    8'h21: p11 <= 8'hfd;
    8'h22: p11 <= 8'h93;
    8'h23: p11 <= 8'h26;
    8'h24: p11 <= 8'h36;
    8'h25: p11 <= 8'h3f;
    8'h26: p11 <= 8'hf7;
    8'h27: p11 <= 8'hcc;
    8'h28: p11 <= 8'h34;
    8'h29: p11 <= 8'ha5;
    8'h2a: p11 <= 8'he5;
    8'h2b: p11 <= 8'hf1;
    8'h2c: p11 <= 8'h71;
    8'h2d: p11 <= 8'hd8;
    8'h2e: p11 <= 8'h31;
    8'h2f: p11 <= 8'h15;
    8'h30: p11 <= 8'h04;
    8'h31: p11 <= 8'hc7;
    8'h32: p11 <= 8'h23;
    8'h33: p11 <= 8'hc3;
    8'h34: p11 <= 8'h18;
    8'h35: p11 <= 8'h96;
    8'h36: p11 <= 8'h05;
    8'h37: p11 <= 8'h9a;
    8'h38: p11 <= 8'h07;
    8'h39: p11 <= 8'h12;
    8'h3a: p11 <= 8'h80;
    8'h3b: p11 <= 8'he2;
    8'h3c: p11 <= 8'heb;
    8'h3d: p11 <= 8'h27;
    8'h3e: p11 <= 8'hb2;
    8'h3f: p11 <= 8'h75;
    8'h40: p11 <= 8'h09;
    8'h41: p11 <= 8'h83;
    8'h42: p11 <= 8'h2c;
    8'h43: p11 <= 8'h1a;
    8'h44: p11 <= 8'h1b;
    8'h45: p11 <= 8'h6e;
    8'h46: p11 <= 8'h5a;
    8'h47: p11 <= 8'ha0;
    8'h48: p11 <= 8'h52;
    8'h49: p11 <= 8'h3b;
    8'h4a: p11 <= 8'hd6;
    8'h4b: p11 <= 8'hb3;
    8'h4c: p11 <= 8'h29;
    8'h4d: p11 <= 8'he3;
    8'h4e: p11 <= 8'h2f;
    8'h4f: p11 <= 8'h84;
    8'h50: p11 <= 8'h53;
    8'h51: p11 <= 8'hd1;
    8'h52: p11 <= 8'h00;
    8'h53: p11 <= 8'hed;
    8'h54: p11 <= 8'h20;
    8'h55: p11 <= 8'hfc;
    8'h56: p11 <= 8'hb1;
    8'h57: p11 <= 8'h5b;
    8'h58: p11 <= 8'h6a;
    8'h59: p11 <= 8'hcb;
    8'h5a: p11 <= 8'hbe;
    8'h5b: p11 <= 8'h39;
    8'h5c: p11 <= 8'h4a;
    8'h5d: p11 <= 8'h4c;
    8'h5e: p11 <= 8'h58;
    8'h5f: p11 <= 8'hcf;
    8'h60: p11 <= 8'hd0;
    8'h61: p11 <= 8'hef;
    8'h62: p11 <= 8'haa;
    8'h63: p11 <= 8'hfb;
    8'h64: p11 <= 8'h43;
    8'h65: p11 <= 8'h4d;
    8'h66: p11 <= 8'h33;
    8'h67: p11 <= 8'h85;
    8'h68: p11 <= 8'h45;
    8'h69: p11 <= 8'hf9;
    8'h6a: p11 <= 8'h02;
    8'h6b: p11 <= 8'h7f;
    8'h6c: p11 <= 8'h50;
    8'h6d: p11 <= 8'h3c;
    8'h6e: p11 <= 8'h9f;
    8'h6f: p11 <= 8'ha8;
    8'h70: p11 <= 8'h51;
    8'h71: p11 <= 8'ha3;
    8'h72: p11 <= 8'h40;
    8'h73: p11 <= 8'h8f;
    8'h74: p11 <= 8'h92;
    8'h75: p11 <= 8'h9d;
    8'h76: p11 <= 8'h38;
    8'h77: p11 <= 8'hf5;
    8'h78: p11 <= 8'hbc;
    8'h79: p11 <= 8'hb6;
    8'h7a: p11 <= 8'hda;
    8'h7b: p11 <= 8'h21;
    8'h7c: p11 <= 8'h10;
    8'h7d: p11 <= 8'hff;
    8'h7e: p11 <= 8'hf3;
    8'h7f: p11 <= 8'hd2;
    8'h80: p11 <= 8'hcd;
    8'h81: p11 <= 8'h0c;
    8'h82: p11 <= 8'h13;
    8'h83: p11 <= 8'hec;
    8'h84: p11 <= 8'h5f;
    8'h85: p11 <= 8'h97;
    8'h86: p11 <= 8'h44;
    8'h87: p11 <= 8'h17;
    8'h88: p11 <= 8'hc4;
    8'h89: p11 <= 8'ha7;
    8'h8a: p11 <= 8'h7e;
    8'h8b: p11 <= 8'h3d;
    8'h8c: p11 <= 8'h64;
    8'h8d: p11 <= 8'h5d;
    8'h8e: p11 <= 8'h19;
    8'h8f: p11 <= 8'h73;
    8'h90: p11 <= 8'h60;
    8'h91: p11 <= 8'h81;
    8'h92: p11 <= 8'h4f;
    8'h93: p11 <= 8'hdc;
    8'h94: p11 <= 8'h22;
    8'h95: p11 <= 8'h2a;
    8'h96: p11 <= 8'h90;
    8'h97: p11 <= 8'h88;
    8'h98: p11 <= 8'h46;
    8'h99: p11 <= 8'hee;
    8'h9a: p11 <= 8'hb8;
    8'h9b: p11 <= 8'h14;
    8'h9c: p11 <= 8'hde;
    8'h9d: p11 <= 8'h5e;
    8'h9e: p11 <= 8'h0b;
    8'h9f: p11 <= 8'hdb;
    8'ha0: p11 <= 8'he0;
    8'ha1: p11 <= 8'h32;
    8'ha2: p11 <= 8'h3a;
    8'ha3: p11 <= 8'h0a;
    8'ha4: p11 <= 8'h49;
    8'ha5: p11 <= 8'h06;
    8'ha6: p11 <= 8'h24;
    8'ha7: p11 <= 8'h5c;
    8'ha8: p11 <= 8'hc2;
    8'ha9: p11 <= 8'hd3;
    8'haa: p11 <= 8'hac;
    8'hab: p11 <= 8'h62;
    8'hac: p11 <= 8'h91;
    8'had: p11 <= 8'h95;
    8'hae: p11 <= 8'he4;
    8'haf: p11 <= 8'h79;
    8'hb0: p11 <= 8'he7;
    8'hb1: p11 <= 8'hc8;
    8'hb2: p11 <= 8'h37;
    8'hb3: p11 <= 8'h6d;
    8'hb4: p11 <= 8'h8d;
    8'hb5: p11 <= 8'hd5;
    8'hb6: p11 <= 8'h4e;
    8'hb7: p11 <= 8'ha9;
    8'hb8: p11 <= 8'h6c;
    8'hb9: p11 <= 8'h56;
    8'hba: p11 <= 8'hf4;
    8'hbb: p11 <= 8'hea;
    8'hbc: p11 <= 8'h65;
    8'hbd: p11 <= 8'h7a;
    8'hbe: p11 <= 8'hae;
    8'hbf: p11 <= 8'h08;
    8'hc0: p11 <= 8'hba;
    8'hc1: p11 <= 8'h78;
    8'hc2: p11 <= 8'h25;
    8'hc3: p11 <= 8'h2e;
    8'hc4: p11 <= 8'h1c;
    8'hc5: p11 <= 8'ha6;
    8'hc6: p11 <= 8'hb4;
    8'hc7: p11 <= 8'hc6;
    8'hc8: p11 <= 8'he8;
    8'hc9: p11 <= 8'hdd;
    8'hca: p11 <= 8'h74;
    8'hcb: p11 <= 8'h1f;
    8'hcc: p11 <= 8'h4b;
    8'hcd: p11 <= 8'hbd;
    8'hce: p11 <= 8'h8b;
    8'hcf: p11 <= 8'h8a;
    8'hd0: p11 <= 8'h70;
    8'hd1: p11 <= 8'h3e;
    8'hd2: p11 <= 8'hb5;
    8'hd3: p11 <= 8'h66;
    8'hd4: p11 <= 8'h48;
    8'hd5: p11 <= 8'h03;
    8'hd6: p11 <= 8'hf6;
    8'hd7: p11 <= 8'h0e;
    8'hd8: p11 <= 8'h61;
    8'hd9: p11 <= 8'h35;
    8'hda: p11 <= 8'h57;
    8'hdb: p11 <= 8'hb9;
    8'hdc: p11 <= 8'h86;
    8'hdd: p11 <= 8'hc1;
    8'hde: p11 <= 8'h1d;
    8'hdf: p11 <= 8'h9e;
    8'he0: p11 <= 8'he1;
    8'he1: p11 <= 8'hf8;
    8'he2: p11 <= 8'h98;
    8'he3: p11 <= 8'h11;
    8'he4: p11 <= 8'h69;
    8'he5: p11 <= 8'hd9;
    8'he6: p11 <= 8'h8e;
    8'he7: p11 <= 8'h94;
    8'he8: p11 <= 8'h9b;
    8'he9: p11 <= 8'h1e;
    8'hea: p11 <= 8'h87;
    8'heb: p11 <= 8'he9;
    8'hec: p11 <= 8'hce;
    8'hed: p11 <= 8'h55;
    8'hee: p11 <= 8'h28;
    8'hef: p11 <= 8'hdf;
    8'hf0: p11 <= 8'h8c;
    8'hf1: p11 <= 8'ha1;
    8'hf2: p11 <= 8'h89;
    8'hf3: p11 <= 8'h0d;
    8'hf4: p11 <= 8'hbf;
    8'hf5: p11 <= 8'he6;
    8'hf6: p11 <= 8'h42;
    8'hf7: p11 <= 8'h68;
    8'hf8: p11 <= 8'h41;
    8'hf9: p11 <= 8'h99;
    8'hfa: p11 <= 8'h2d;
    8'hfb: p11 <= 8'h0f;
    8'hfc: p11 <= 8'hb0;
    8'hfd: p11 <= 8'h54;
    8'hfe: p11 <= 8'hbb;
    8'hff: p11 <= 8'h16;
    endcase
	
    // Third Portion
    case (s1[23:16])
    8'h00: p12 <= 8'h63;
    8'h01: p12 <= 8'h7c;
    8'h02: p12 <= 8'h77;
    8'h03: p12 <= 8'h7b;
    8'h04: p12 <= 8'hf2;
    8'h05: p12 <= 8'h6b;
    8'h06: p12 <= 8'h6f;
    8'h07: p12 <= 8'hc5;
    8'h08: p12 <= 8'h30;
    8'h09: p12 <= 8'h01;
    8'h0a: p12 <= 8'h67;
    8'h0b: p12 <= 8'h2b;
    8'h0c: p12 <= 8'hfe;
    8'h0d: p12 <= 8'hd7;
    8'h0e: p12 <= 8'hab;
    8'h0f: p12 <= 8'h76;
    8'h10: p12 <= 8'hca;
    8'h11: p12 <= 8'h82;
    8'h12: p12 <= 8'hc9;
    8'h13: p12 <= 8'h7d;
    8'h14: p12 <= 8'hfa;
    8'h15: p12 <= 8'h59;
    8'h16: p12 <= 8'h47;
    8'h17: p12 <= 8'hf0;
    8'h18: p12 <= 8'had;
    8'h19: p12 <= 8'hd4;
    8'h1a: p12 <= 8'ha2;
    8'h1b: p12 <= 8'haf;
    8'h1c: p12 <= 8'h9c;
    8'h1d: p12 <= 8'ha4;
    8'h1e: p12 <= 8'h72;
    8'h1f: p12 <= 8'hc0;
    8'h20: p12 <= 8'hb7;
    8'h21: p12 <= 8'hfd;
    8'h22: p12 <= 8'h93;
    8'h23: p12 <= 8'h26;
    8'h24: p12 <= 8'h36;
    8'h25: p12 <= 8'h3f;
    8'h26: p12 <= 8'hf7;
    8'h27: p12 <= 8'hcc;
    8'h28: p12 <= 8'h34;
    8'h29: p12 <= 8'ha5;
    8'h2a: p12 <= 8'he5;
    8'h2b: p12 <= 8'hf1;
    8'h2c: p12 <= 8'h71;
    8'h2d: p12 <= 8'hd8;
    8'h2e: p12 <= 8'h31;
    8'h2f: p12 <= 8'h15;
    8'h30: p12 <= 8'h04;
    8'h31: p12 <= 8'hc7;
    8'h32: p12 <= 8'h23;
    8'h33: p12 <= 8'hc3;
    8'h34: p12 <= 8'h18;
    8'h35: p12 <= 8'h96;
    8'h36: p12 <= 8'h05;
    8'h37: p12 <= 8'h9a;
    8'h38: p12 <= 8'h07;
    8'h39: p12 <= 8'h12;
    8'h3a: p12 <= 8'h80;
    8'h3b: p12 <= 8'he2;
    8'h3c: p12 <= 8'heb;
    8'h3d: p12 <= 8'h27;
    8'h3e: p12 <= 8'hb2;
    8'h3f: p12 <= 8'h75;
    8'h40: p12 <= 8'h09;
    8'h41: p12 <= 8'h83;
    8'h42: p12 <= 8'h2c;
    8'h43: p12 <= 8'h1a;
    8'h44: p12 <= 8'h1b;
    8'h45: p12 <= 8'h6e;
    8'h46: p12 <= 8'h5a;
    8'h47: p12 <= 8'ha0;
    8'h48: p12 <= 8'h52;
    8'h49: p12 <= 8'h3b;
    8'h4a: p12 <= 8'hd6;
    8'h4b: p12 <= 8'hb3;
    8'h4c: p12 <= 8'h29;
    8'h4d: p12 <= 8'he3;
    8'h4e: p12 <= 8'h2f;
    8'h4f: p12 <= 8'h84;
    8'h50: p12 <= 8'h53;
    8'h51: p12 <= 8'hd1;
    8'h52: p12 <= 8'h00;
    8'h53: p12 <= 8'hed;
    8'h54: p12 <= 8'h20;
    8'h55: p12 <= 8'hfc;
    8'h56: p12 <= 8'hb1;
    8'h57: p12 <= 8'h5b;
    8'h58: p12 <= 8'h6a;
    8'h59: p12 <= 8'hcb;
    8'h5a: p12 <= 8'hbe;
    8'h5b: p12 <= 8'h39;
    8'h5c: p12 <= 8'h4a;
    8'h5d: p12 <= 8'h4c;
    8'h5e: p12 <= 8'h58;
    8'h5f: p12 <= 8'hcf;
    8'h60: p12 <= 8'hd0;
    8'h61: p12 <= 8'hef;
    8'h62: p12 <= 8'haa;
    8'h63: p12 <= 8'hfb;
    8'h64: p12 <= 8'h43;
    8'h65: p12 <= 8'h4d;
    8'h66: p12 <= 8'h33;
    8'h67: p12 <= 8'h85;
    8'h68: p12 <= 8'h45;
    8'h69: p12 <= 8'hf9;
    8'h6a: p12 <= 8'h02;
    8'h6b: p12 <= 8'h7f;
    8'h6c: p12 <= 8'h50;
    8'h6d: p12 <= 8'h3c;
    8'h6e: p12 <= 8'h9f;
    8'h6f: p12 <= 8'ha8;
    8'h70: p12 <= 8'h51;
    8'h71: p12 <= 8'ha3;
    8'h72: p12 <= 8'h40;
    8'h73: p12 <= 8'h8f;
    8'h74: p12 <= 8'h92;
    8'h75: p12 <= 8'h9d;
    8'h76: p12 <= 8'h38;
    8'h77: p12 <= 8'hf5;
    8'h78: p12 <= 8'hbc;
    8'h79: p12 <= 8'hb6;
    8'h7a: p12 <= 8'hda;
    8'h7b: p12 <= 8'h21;
    8'h7c: p12 <= 8'h10;
    8'h7d: p12 <= 8'hff;
    8'h7e: p12 <= 8'hf3;
    8'h7f: p12 <= 8'hd2;
    8'h80: p12 <= 8'hcd;
    8'h81: p12 <= 8'h0c;
    8'h82: p12 <= 8'h13;
    8'h83: p12 <= 8'hec;
    8'h84: p12 <= 8'h5f;
    8'h85: p12 <= 8'h97;
    8'h86: p12 <= 8'h44;
    8'h87: p12 <= 8'h17;
    8'h88: p12 <= 8'hc4;
    8'h89: p12 <= 8'ha7;
    8'h8a: p12 <= 8'h7e;
    8'h8b: p12 <= 8'h3d;
    8'h8c: p12 <= 8'h64;
    8'h8d: p12 <= 8'h5d;
    8'h8e: p12 <= 8'h19;
    8'h8f: p12 <= 8'h73;
    8'h90: p12 <= 8'h60;
    8'h91: p12 <= 8'h81;
    8'h92: p12 <= 8'h4f;
    8'h93: p12 <= 8'hdc;
    8'h94: p12 <= 8'h22;
    8'h95: p12 <= 8'h2a;
    8'h96: p12 <= 8'h90;
    8'h97: p12 <= 8'h88;
    8'h98: p12 <= 8'h46;
    8'h99: p12 <= 8'hee;
    8'h9a: p12 <= 8'hb8;
    8'h9b: p12 <= 8'h14;
    8'h9c: p12 <= 8'hde;
    8'h9d: p12 <= 8'h5e;
    8'h9e: p12 <= 8'h0b;
    8'h9f: p12 <= 8'hdb;
    8'ha0: p12 <= 8'he0;
    8'ha1: p12 <= 8'h32;
    8'ha2: p12 <= 8'h3a;
    8'ha3: p12 <= 8'h0a;
    8'ha4: p12 <= 8'h49;
    8'ha5: p12 <= 8'h06;
    8'ha6: p12 <= 8'h24;
    8'ha7: p12 <= 8'h5c;
    8'ha8: p12 <= 8'hc2;
    8'ha9: p12 <= 8'hd3;
    8'haa: p12 <= 8'hac;
    8'hab: p12 <= 8'h62;
    8'hac: p12 <= 8'h91;
    8'had: p12 <= 8'h95;
    8'hae: p12 <= 8'he4;
    8'haf: p12 <= 8'h79;
    8'hb0: p12 <= 8'he7;
    8'hb1: p12 <= 8'hc8;
    8'hb2: p12 <= 8'h37;
    8'hb3: p12 <= 8'h6d;
    8'hb4: p12 <= 8'h8d;
    8'hb5: p12 <= 8'hd5;
    8'hb6: p12 <= 8'h4e;
    8'hb7: p12 <= 8'ha9;
    8'hb8: p12 <= 8'h6c;
    8'hb9: p12 <= 8'h56;
    8'hba: p12 <= 8'hf4;
    8'hbb: p12 <= 8'hea;
    8'hbc: p12 <= 8'h65;
    8'hbd: p12 <= 8'h7a;
    8'hbe: p12 <= 8'hae;
    8'hbf: p12 <= 8'h08;
    8'hc0: p12 <= 8'hba;
    8'hc1: p12 <= 8'h78;
    8'hc2: p12 <= 8'h25;
    8'hc3: p12 <= 8'h2e;
    8'hc4: p12 <= 8'h1c;
    8'hc5: p12 <= 8'ha6;
    8'hc6: p12 <= 8'hb4;
    8'hc7: p12 <= 8'hc6;
    8'hc8: p12 <= 8'he8;
    8'hc9: p12 <= 8'hdd;
    8'hca: p12 <= 8'h74;
    8'hcb: p12 <= 8'h1f;
    8'hcc: p12 <= 8'h4b;
    8'hcd: p12 <= 8'hbd;
    8'hce: p12 <= 8'h8b;
    8'hcf: p12 <= 8'h8a;
    8'hd0: p12 <= 8'h70;
    8'hd1: p12 <= 8'h3e;
    8'hd2: p12 <= 8'hb5;
    8'hd3: p12 <= 8'h66;
    8'hd4: p12 <= 8'h48;
    8'hd5: p12 <= 8'h03;
    8'hd6: p12 <= 8'hf6;
    8'hd7: p12 <= 8'h0e;
    8'hd8: p12 <= 8'h61;
    8'hd9: p12 <= 8'h35;
    8'hda: p12 <= 8'h57;
    8'hdb: p12 <= 8'hb9;
    8'hdc: p12 <= 8'h86;
    8'hdd: p12 <= 8'hc1;
    8'hde: p12 <= 8'h1d;
    8'hdf: p12 <= 8'h9e;
    8'he0: p12 <= 8'he1;
    8'he1: p12 <= 8'hf8;
    8'he2: p12 <= 8'h98;
    8'he3: p12 <= 8'h11;
    8'he4: p12 <= 8'h69;
    8'he5: p12 <= 8'hd9;
    8'he6: p12 <= 8'h8e;
    8'he7: p12 <= 8'h94;
    8'he8: p12 <= 8'h9b;
    8'he9: p12 <= 8'h1e;
    8'hea: p12 <= 8'h87;
    8'heb: p12 <= 8'he9;
    8'hec: p12 <= 8'hce;
    8'hed: p12 <= 8'h55;
    8'hee: p12 <= 8'h28;
    8'hef: p12 <= 8'hdf;
    8'hf0: p12 <= 8'h8c;
    8'hf1: p12 <= 8'ha1;
    8'hf2: p12 <= 8'h89;
    8'hf3: p12 <= 8'h0d;
    8'hf4: p12 <= 8'hbf;
    8'hf5: p12 <= 8'he6;
    8'hf6: p12 <= 8'h42;
    8'hf7: p12 <= 8'h68;
    8'hf8: p12 <= 8'h41;
    8'hf9: p12 <= 8'h99;
    8'hfa: p12 <= 8'h2d;
    8'hfb: p12 <= 8'h0f;
    8'hfc: p12 <= 8'hb0;
    8'hfd: p12 <= 8'h54;
    8'hfe: p12 <= 8'hbb;
    8'hff: p12 <= 8'h16;
    endcase
	
    // Fourth Portion
    case (s1[31:24])
    8'h00: p13 <= 8'h63;
    8'h01: p13 <= 8'h7c;
    8'h02: p13 <= 8'h77;
    8'h03: p13 <= 8'h7b;
    8'h04: p13 <= 8'hf2;
    8'h05: p13 <= 8'h6b;
    8'h06: p13 <= 8'h6f;
    8'h07: p13 <= 8'hc5;
    8'h08: p13 <= 8'h30;
    8'h09: p13 <= 8'h01;
    8'h0a: p13 <= 8'h67;
    8'h0b: p13 <= 8'h2b;
    8'h0c: p13 <= 8'hfe;
    8'h0d: p13 <= 8'hd7;
    8'h0e: p13 <= 8'hab;
    8'h0f: p13 <= 8'h76;
    8'h10: p13 <= 8'hca;
    8'h11: p13 <= 8'h82;
    8'h12: p13 <= 8'hc9;
    8'h13: p13 <= 8'h7d;
    8'h14: p13 <= 8'hfa;
    8'h15: p13 <= 8'h59;
    8'h16: p13 <= 8'h47;
    8'h17: p13 <= 8'hf0;
    8'h18: p13 <= 8'had;
    8'h19: p13 <= 8'hd4;
    8'h1a: p13 <= 8'ha2;
    8'h1b: p13 <= 8'haf;
    8'h1c: p13 <= 8'h9c;
    8'h1d: p13 <= 8'ha4;
    8'h1e: p13 <= 8'h72;
    8'h1f: p13 <= 8'hc0;
    8'h20: p13 <= 8'hb7;
    8'h21: p13 <= 8'hfd;
    8'h22: p13 <= 8'h93;
    8'h23: p13 <= 8'h26;
    8'h24: p13 <= 8'h36;
    8'h25: p13 <= 8'h3f;
    8'h26: p13 <= 8'hf7;
    8'h27: p13 <= 8'hcc;
    8'h28: p13 <= 8'h34;
    8'h29: p13 <= 8'ha5;
    8'h2a: p13 <= 8'he5;
    8'h2b: p13 <= 8'hf1;
    8'h2c: p13 <= 8'h71;
    8'h2d: p13 <= 8'hd8;
    8'h2e: p13 <= 8'h31;
    8'h2f: p13 <= 8'h15;
    8'h30: p13 <= 8'h04;
    8'h31: p13 <= 8'hc7;
    8'h32: p13 <= 8'h23;
    8'h33: p13 <= 8'hc3;
    8'h34: p13 <= 8'h18;
    8'h35: p13 <= 8'h96;
    8'h36: p13 <= 8'h05;
    8'h37: p13 <= 8'h9a;
    8'h38: p13 <= 8'h07;
    8'h39: p13 <= 8'h12;
    8'h3a: p13 <= 8'h80;
    8'h3b: p13 <= 8'he2;
    8'h3c: p13 <= 8'heb;
    8'h3d: p13 <= 8'h27;
    8'h3e: p13 <= 8'hb2;
    8'h3f: p13 <= 8'h75;
    8'h40: p13 <= 8'h09;
    8'h41: p13 <= 8'h83;
    8'h42: p13 <= 8'h2c;
    8'h43: p13 <= 8'h1a;
    8'h44: p13 <= 8'h1b;
    8'h45: p13 <= 8'h6e;
    8'h46: p13 <= 8'h5a;
    8'h47: p13 <= 8'ha0;
    8'h48: p13 <= 8'h52;
    8'h49: p13 <= 8'h3b;
    8'h4a: p13 <= 8'hd6;
    8'h4b: p13 <= 8'hb3;
    8'h4c: p13 <= 8'h29;
    8'h4d: p13 <= 8'he3;
    8'h4e: p13 <= 8'h2f;
    8'h4f: p13 <= 8'h84;
    8'h50: p13 <= 8'h53;
    8'h51: p13 <= 8'hd1;
    8'h52: p13 <= 8'h00;
    8'h53: p13 <= 8'hed;
    8'h54: p13 <= 8'h20;
    8'h55: p13 <= 8'hfc;
    8'h56: p13 <= 8'hb1;
    8'h57: p13 <= 8'h5b;
    8'h58: p13 <= 8'h6a;
    8'h59: p13 <= 8'hcb;
    8'h5a: p13 <= 8'hbe;
    8'h5b: p13 <= 8'h39;
    8'h5c: p13 <= 8'h4a;
    8'h5d: p13 <= 8'h4c;
    8'h5e: p13 <= 8'h58;
    8'h5f: p13 <= 8'hcf;
    8'h60: p13 <= 8'hd0;
    8'h61: p13 <= 8'hef;
    8'h62: p13 <= 8'haa;
    8'h63: p13 <= 8'hfb;
    8'h64: p13 <= 8'h43;
    8'h65: p13 <= 8'h4d;
    8'h66: p13 <= 8'h33;
    8'h67: p13 <= 8'h85;
    8'h68: p13 <= 8'h45;
    8'h69: p13 <= 8'hf9;
    8'h6a: p13 <= 8'h02;
    8'h6b: p13 <= 8'h7f;
    8'h6c: p13 <= 8'h50;
    8'h6d: p13 <= 8'h3c;
    8'h6e: p13 <= 8'h9f;
    8'h6f: p13 <= 8'ha8;
    8'h70: p13 <= 8'h51;
    8'h71: p13 <= 8'ha3;
    8'h72: p13 <= 8'h40;
    8'h73: p13 <= 8'h8f;
    8'h74: p13 <= 8'h92;
    8'h75: p13 <= 8'h9d;
    8'h76: p13 <= 8'h38;
    8'h77: p13 <= 8'hf5;
    8'h78: p13 <= 8'hbc;
    8'h79: p13 <= 8'hb6;
    8'h7a: p13 <= 8'hda;
    8'h7b: p13 <= 8'h21;
    8'h7c: p13 <= 8'h10;
    8'h7d: p13 <= 8'hff;
    8'h7e: p13 <= 8'hf3;
    8'h7f: p13 <= 8'hd2;
    8'h80: p13 <= 8'hcd;
    8'h81: p13 <= 8'h0c;
    8'h82: p13 <= 8'h13;
    8'h83: p13 <= 8'hec;
    8'h84: p13 <= 8'h5f;
    8'h85: p13 <= 8'h97;
    8'h86: p13 <= 8'h44;
    8'h87: p13 <= 8'h17;
    8'h88: p13 <= 8'hc4;
    8'h89: p13 <= 8'ha7;
    8'h8a: p13 <= 8'h7e;
    8'h8b: p13 <= 8'h3d;
    8'h8c: p13 <= 8'h64;
    8'h8d: p13 <= 8'h5d;
    8'h8e: p13 <= 8'h19;
    8'h8f: p13 <= 8'h73;
    8'h90: p13 <= 8'h60;
    8'h91: p13 <= 8'h81;
    8'h92: p13 <= 8'h4f;
    8'h93: p13 <= 8'hdc;
    8'h94: p13 <= 8'h22;
    8'h95: p13 <= 8'h2a;
    8'h96: p13 <= 8'h90;
    8'h97: p13 <= 8'h88;
    8'h98: p13 <= 8'h46;
    8'h99: p13 <= 8'hee;
    8'h9a: p13 <= 8'hb8;
    8'h9b: p13 <= 8'h14;
    8'h9c: p13 <= 8'hde;
    8'h9d: p13 <= 8'h5e;
    8'h9e: p13 <= 8'h0b;
    8'h9f: p13 <= 8'hdb;
    8'ha0: p13 <= 8'he0;
    8'ha1: p13 <= 8'h32;
    8'ha2: p13 <= 8'h3a;
    8'ha3: p13 <= 8'h0a;
    8'ha4: p13 <= 8'h49;
    8'ha5: p13 <= 8'h06;
    8'ha6: p13 <= 8'h24;
    8'ha7: p13 <= 8'h5c;
    8'ha8: p13 <= 8'hc2;
    8'ha9: p13 <= 8'hd3;
    8'haa: p13 <= 8'hac;
    8'hab: p13 <= 8'h62;
    8'hac: p13 <= 8'h91;
    8'had: p13 <= 8'h95;
    8'hae: p13 <= 8'he4;
    8'haf: p13 <= 8'h79;
    8'hb0: p13 <= 8'he7;
    8'hb1: p13 <= 8'hc8;
    8'hb2: p13 <= 8'h37;
    8'hb3: p13 <= 8'h6d;
    8'hb4: p13 <= 8'h8d;
    8'hb5: p13 <= 8'hd5;
    8'hb6: p13 <= 8'h4e;
    8'hb7: p13 <= 8'ha9;
    8'hb8: p13 <= 8'h6c;
    8'hb9: p13 <= 8'h56;
    8'hba: p13 <= 8'hf4;
    8'hbb: p13 <= 8'hea;
    8'hbc: p13 <= 8'h65;
    8'hbd: p13 <= 8'h7a;
    8'hbe: p13 <= 8'hae;
    8'hbf: p13 <= 8'h08;
    8'hc0: p13 <= 8'hba;
    8'hc1: p13 <= 8'h78;
    8'hc2: p13 <= 8'h25;
    8'hc3: p13 <= 8'h2e;
    8'hc4: p13 <= 8'h1c;
    8'hc5: p13 <= 8'ha6;
    8'hc6: p13 <= 8'hb4;
    8'hc7: p13 <= 8'hc6;
    8'hc8: p13 <= 8'he8;
    8'hc9: p13 <= 8'hdd;
    8'hca: p13 <= 8'h74;
    8'hcb: p13 <= 8'h1f;
    8'hcc: p13 <= 8'h4b;
    8'hcd: p13 <= 8'hbd;
    8'hce: p13 <= 8'h8b;
    8'hcf: p13 <= 8'h8a;
    8'hd0: p13 <= 8'h70;
    8'hd1: p13 <= 8'h3e;
    8'hd2: p13 <= 8'hb5;
    8'hd3: p13 <= 8'h66;
    8'hd4: p13 <= 8'h48;
    8'hd5: p13 <= 8'h03;
    8'hd6: p13 <= 8'hf6;
    8'hd7: p13 <= 8'h0e;
    8'hd8: p13 <= 8'h61;
    8'hd9: p13 <= 8'h35;
    8'hda: p13 <= 8'h57;
    8'hdb: p13 <= 8'hb9;
    8'hdc: p13 <= 8'h86;
    8'hdd: p13 <= 8'hc1;
    8'hde: p13 <= 8'h1d;
    8'hdf: p13 <= 8'h9e;
    8'he0: p13 <= 8'he1;
    8'he1: p13 <= 8'hf8;
    8'he2: p13 <= 8'h98;
    8'he3: p13 <= 8'h11;
    8'he4: p13 <= 8'h69;
    8'he5: p13 <= 8'hd9;
    8'he6: p13 <= 8'h8e;
    8'he7: p13 <= 8'h94;
    8'he8: p13 <= 8'h9b;
    8'he9: p13 <= 8'h1e;
    8'hea: p13 <= 8'h87;
    8'heb: p13 <= 8'he9;
    8'hec: p13 <= 8'hce;
    8'hed: p13 <= 8'h55;
    8'hee: p13 <= 8'h28;
    8'hef: p13 <= 8'hdf;
    8'hf0: p13 <= 8'h8c;
    8'hf1: p13 <= 8'ha1;
    8'hf2: p13 <= 8'h89;
    8'hf3: p13 <= 8'h0d;
    8'hf4: p13 <= 8'hbf;
    8'hf5: p13 <= 8'he6;
    8'hf6: p13 <= 8'h42;
    8'hf7: p13 <= 8'h68;
    8'hf8: p13 <= 8'h41;
    8'hf9: p13 <= 8'h99;
    8'hfa: p13 <= 8'h2d;
    8'hfb: p13 <= 8'h0f;
    8'hfc: p13 <= 8'hb0;
    8'hfd: p13 <= 8'h54;
    8'hfe: p13 <= 8'hbb;
    8'hff: p13 <= 8'h16;
    endcase
	
	// **************************** PART S2 ****************************
	
    // First Portion
    case (s2[7:0])
    8'h00: p20 <= 8'h63;
    8'h01: p20 <= 8'h7c;
    8'h02: p20 <= 8'h77;
    8'h03: p20 <= 8'h7b;
    8'h04: p20 <= 8'hf2;
    8'h05: p20 <= 8'h6b;
    8'h06: p20 <= 8'h6f;
    8'h07: p20 <= 8'hc5;
    8'h08: p20 <= 8'h30;
    8'h09: p20 <= 8'h01;
    8'h0a: p20 <= 8'h67;
    8'h0b: p20 <= 8'h2b;
    8'h0c: p20 <= 8'hfe;
    8'h0d: p20 <= 8'hd7;
    8'h0e: p20 <= 8'hab;
    8'h0f: p20 <= 8'h76;
    8'h10: p20 <= 8'hca;
    8'h11: p20 <= 8'h82;
    8'h12: p20 <= 8'hc9;
    8'h13: p20 <= 8'h7d;
    8'h14: p20 <= 8'hfa;
    8'h15: p20 <= 8'h59;
    8'h16: p20 <= 8'h47;
    8'h17: p20 <= 8'hf0;
    8'h18: p20 <= 8'had;
    8'h19: p20 <= 8'hd4;
    8'h1a: p20 <= 8'ha2;
    8'h1b: p20 <= 8'haf;
    8'h1c: p20 <= 8'h9c;
    8'h1d: p20 <= 8'ha4;
    8'h1e: p20 <= 8'h72;
    8'h1f: p20 <= 8'hc0;
    8'h20: p20 <= 8'hb7;
    8'h21: p20 <= 8'hfd;
    8'h22: p20 <= 8'h93;
    8'h23: p20 <= 8'h26;
    8'h24: p20 <= 8'h36;
    8'h25: p20 <= 8'h3f;
    8'h26: p20 <= 8'hf7;
    8'h27: p20 <= 8'hcc;
    8'h28: p20 <= 8'h34;
    8'h29: p20 <= 8'ha5;
    8'h2a: p20 <= 8'he5;
    8'h2b: p20 <= 8'hf1;
    8'h2c: p20 <= 8'h71;
    8'h2d: p20 <= 8'hd8;
    8'h2e: p20 <= 8'h31;
    8'h2f: p20 <= 8'h15;
    8'h30: p20 <= 8'h04;
    8'h31: p20 <= 8'hc7;
    8'h32: p20 <= 8'h23;
    8'h33: p20 <= 8'hc3;
    8'h34: p20 <= 8'h18;
    8'h35: p20 <= 8'h96;
    8'h36: p20 <= 8'h05;
    8'h37: p20 <= 8'h9a;
    8'h38: p20 <= 8'h07;
    8'h39: p20 <= 8'h12;
    8'h3a: p20 <= 8'h80;
    8'h3b: p20 <= 8'he2;
    8'h3c: p20 <= 8'heb;
    8'h3d: p20 <= 8'h27;
    8'h3e: p20 <= 8'hb2;
    8'h3f: p20 <= 8'h75;
    8'h40: p20 <= 8'h09;
    8'h41: p20 <= 8'h83;
    8'h42: p20 <= 8'h2c;
    8'h43: p20 <= 8'h1a;
    8'h44: p20 <= 8'h1b;
    8'h45: p20 <= 8'h6e;
    8'h46: p20 <= 8'h5a;
    8'h47: p20 <= 8'ha0;
    8'h48: p20 <= 8'h52;
    8'h49: p20 <= 8'h3b;
    8'h4a: p20 <= 8'hd6;
    8'h4b: p20 <= 8'hb3;
    8'h4c: p20 <= 8'h29;
    8'h4d: p20 <= 8'he3;
    8'h4e: p20 <= 8'h2f;
    8'h4f: p20 <= 8'h84;
    8'h50: p20 <= 8'h53;
    8'h51: p20 <= 8'hd1;
    8'h52: p20 <= 8'h00;
    8'h53: p20 <= 8'hed;
    8'h54: p20 <= 8'h20;
    8'h55: p20 <= 8'hfc;
    8'h56: p20 <= 8'hb1;
    8'h57: p20 <= 8'h5b;
    8'h58: p20 <= 8'h6a;
    8'h59: p20 <= 8'hcb;
    8'h5a: p20 <= 8'hbe;
    8'h5b: p20 <= 8'h39;
    8'h5c: p20 <= 8'h4a;
    8'h5d: p20 <= 8'h4c;
    8'h5e: p20 <= 8'h58;
    8'h5f: p20 <= 8'hcf;
    8'h60: p20 <= 8'hd0;
    8'h61: p20 <= 8'hef;
    8'h62: p20 <= 8'haa;
    8'h63: p20 <= 8'hfb;
    8'h64: p20 <= 8'h43;
    8'h65: p20 <= 8'h4d;
    8'h66: p20 <= 8'h33;
    8'h67: p20 <= 8'h85;
    8'h68: p20 <= 8'h45;
    8'h69: p20 <= 8'hf9;
    8'h6a: p20 <= 8'h02;
    8'h6b: p20 <= 8'h7f;
    8'h6c: p20 <= 8'h50;
    8'h6d: p20 <= 8'h3c;
    8'h6e: p20 <= 8'h9f;
    8'h6f: p20 <= 8'ha8;
    8'h70: p20 <= 8'h51;
    8'h71: p20 <= 8'ha3;
    8'h72: p20 <= 8'h40;
    8'h73: p20 <= 8'h8f;
    8'h74: p20 <= 8'h92;
    8'h75: p20 <= 8'h9d;
    8'h76: p20 <= 8'h38;
    8'h77: p20 <= 8'hf5;
    8'h78: p20 <= 8'hbc;
    8'h79: p20 <= 8'hb6;
    8'h7a: p20 <= 8'hda;
    8'h7b: p20 <= 8'h21;
    8'h7c: p20 <= 8'h10;
    8'h7d: p20 <= 8'hff;
    8'h7e: p20 <= 8'hf3;
    8'h7f: p20 <= 8'hd2;
    8'h80: p20 <= 8'hcd;
    8'h81: p20 <= 8'h0c;
    8'h82: p20 <= 8'h13;
    8'h83: p20 <= 8'hec;
    8'h84: p20 <= 8'h5f;
    8'h85: p20 <= 8'h97;
    8'h86: p20 <= 8'h44;
    8'h87: p20 <= 8'h17;
    8'h88: p20 <= 8'hc4;
    8'h89: p20 <= 8'ha7;
    8'h8a: p20 <= 8'h7e;
    8'h8b: p20 <= 8'h3d;
    8'h8c: p20 <= 8'h64;
    8'h8d: p20 <= 8'h5d;
    8'h8e: p20 <= 8'h19;
    8'h8f: p20 <= 8'h73;
    8'h90: p20 <= 8'h60;
    8'h91: p20 <= 8'h81;
    8'h92: p20 <= 8'h4f;
    8'h93: p20 <= 8'hdc;
    8'h94: p20 <= 8'h22;
    8'h95: p20 <= 8'h2a;
    8'h96: p20 <= 8'h90;
    8'h97: p20 <= 8'h88;
    8'h98: p20 <= 8'h46;
    8'h99: p20 <= 8'hee;
    8'h9a: p20 <= 8'hb8;
    8'h9b: p20 <= 8'h14;
    8'h9c: p20 <= 8'hde;
    8'h9d: p20 <= 8'h5e;
    8'h9e: p20 <= 8'h0b;
    8'h9f: p20 <= 8'hdb;
    8'ha0: p20 <= 8'he0;
    8'ha1: p20 <= 8'h32;
    8'ha2: p20 <= 8'h3a;
    8'ha3: p20 <= 8'h0a;
    8'ha4: p20 <= 8'h49;
    8'ha5: p20 <= 8'h06;
    8'ha6: p20 <= 8'h24;
    8'ha7: p20 <= 8'h5c;
    8'ha8: p20 <= 8'hc2;
    8'ha9: p20 <= 8'hd3;
    8'haa: p20 <= 8'hac;
    8'hab: p20 <= 8'h62;
    8'hac: p20 <= 8'h91;
    8'had: p20 <= 8'h95;
    8'hae: p20 <= 8'he4;
    8'haf: p20 <= 8'h79;
    8'hb0: p20 <= 8'he7;
    8'hb1: p20 <= 8'hc8;
    8'hb2: p20 <= 8'h37;
    8'hb3: p20 <= 8'h6d;
    8'hb4: p20 <= 8'h8d;
    8'hb5: p20 <= 8'hd5;
    8'hb6: p20 <= 8'h4e;
    8'hb7: p20 <= 8'ha9;
    8'hb8: p20 <= 8'h6c;
    8'hb9: p20 <= 8'h56;
    8'hba: p20 <= 8'hf4;
    8'hbb: p20 <= 8'hea;
    8'hbc: p20 <= 8'h65;
    8'hbd: p20 <= 8'h7a;
    8'hbe: p20 <= 8'hae;
    8'hbf: p20 <= 8'h08;
    8'hc0: p20 <= 8'hba;
    8'hc1: p20 <= 8'h78;
    8'hc2: p20 <= 8'h25;
    8'hc3: p20 <= 8'h2e;
    8'hc4: p20 <= 8'h1c;
    8'hc5: p20 <= 8'ha6;
    8'hc6: p20 <= 8'hb4;
    8'hc7: p20 <= 8'hc6;
    8'hc8: p20 <= 8'he8;
    8'hc9: p20 <= 8'hdd;
    8'hca: p20 <= 8'h74;
    8'hcb: p20 <= 8'h1f;
    8'hcc: p20 <= 8'h4b;
    8'hcd: p20 <= 8'hbd;
    8'hce: p20 <= 8'h8b;
    8'hcf: p20 <= 8'h8a;
    8'hd0: p20 <= 8'h70;
    8'hd1: p20 <= 8'h3e;
    8'hd2: p20 <= 8'hb5;
    8'hd3: p20 <= 8'h66;
    8'hd4: p20 <= 8'h48;
    8'hd5: p20 <= 8'h03;
    8'hd6: p20 <= 8'hf6;
    8'hd7: p20 <= 8'h0e;
    8'hd8: p20 <= 8'h61;
    8'hd9: p20 <= 8'h35;
    8'hda: p20 <= 8'h57;
    8'hdb: p20 <= 8'hb9;
    8'hdc: p20 <= 8'h86;
    8'hdd: p20 <= 8'hc1;
    8'hde: p20 <= 8'h1d;
    8'hdf: p20 <= 8'h9e;
    8'he0: p20 <= 8'he1;
    8'he1: p20 <= 8'hf8;
    8'he2: p20 <= 8'h98;
    8'he3: p20 <= 8'h11;
    8'he4: p20 <= 8'h69;
    8'he5: p20 <= 8'hd9;
    8'he6: p20 <= 8'h8e;
    8'he7: p20 <= 8'h94;
    8'he8: p20 <= 8'h9b;
    8'he9: p20 <= 8'h1e;
    8'hea: p20 <= 8'h87;
    8'heb: p20 <= 8'he9;
    8'hec: p20 <= 8'hce;
    8'hed: p20 <= 8'h55;
    8'hee: p20 <= 8'h28;
    8'hef: p20 <= 8'hdf;
    8'hf0: p20 <= 8'h8c;
    8'hf1: p20 <= 8'ha1;
    8'hf2: p20 <= 8'h89;
    8'hf3: p20 <= 8'h0d;
    8'hf4: p20 <= 8'hbf;
    8'hf5: p20 <= 8'he6;
    8'hf6: p20 <= 8'h42;
    8'hf7: p20 <= 8'h68;
    8'hf8: p20 <= 8'h41;
    8'hf9: p20 <= 8'h99;
    8'hfa: p20 <= 8'h2d;
    8'hfb: p20 <= 8'h0f;
    8'hfc: p20 <= 8'hb0;
    8'hfd: p20 <= 8'h54;
    8'hfe: p20 <= 8'hbb;
    8'hff: p20 <= 8'h16;
    endcase
	
    // Second Portion
    case (s2[15:8])
    8'h00: p21 <= 8'h63;
    8'h01: p21 <= 8'h7c;
    8'h02: p21 <= 8'h77;
    8'h03: p21 <= 8'h7b;
    8'h04: p21 <= 8'hf2;
    8'h05: p21 <= 8'h6b;
    8'h06: p21 <= 8'h6f;
    8'h07: p21 <= 8'hc5;
    8'h08: p21 <= 8'h30;
    8'h09: p21 <= 8'h01;
    8'h0a: p21 <= 8'h67;
    8'h0b: p21 <= 8'h2b;
    8'h0c: p21 <= 8'hfe;
    8'h0d: p21 <= 8'hd7;
    8'h0e: p21 <= 8'hab;
    8'h0f: p21 <= 8'h76;
    8'h10: p21 <= 8'hca;
    8'h11: p21 <= 8'h82;
    8'h12: p21 <= 8'hc9;
    8'h13: p21 <= 8'h7d;
    8'h14: p21 <= 8'hfa;
    8'h15: p21 <= 8'h59;
    8'h16: p21 <= 8'h47;
    8'h17: p21 <= 8'hf0;
    8'h18: p21 <= 8'had;
    8'h19: p21 <= 8'hd4;
    8'h1a: p21 <= 8'ha2;
    8'h1b: p21 <= 8'haf;
    8'h1c: p21 <= 8'h9c;
    8'h1d: p21 <= 8'ha4;
    8'h1e: p21 <= 8'h72;
    8'h1f: p21 <= 8'hc0;
    8'h20: p21 <= 8'hb7;
    8'h21: p21 <= 8'hfd;
    8'h22: p21 <= 8'h93;
    8'h23: p21 <= 8'h26;
    8'h24: p21 <= 8'h36;
    8'h25: p21 <= 8'h3f;
    8'h26: p21 <= 8'hf7;
    8'h27: p21 <= 8'hcc;
    8'h28: p21 <= 8'h34;
    8'h29: p21 <= 8'ha5;
    8'h2a: p21 <= 8'he5;
    8'h2b: p21 <= 8'hf1;
    8'h2c: p21 <= 8'h71;
    8'h2d: p21 <= 8'hd8;
    8'h2e: p21 <= 8'h31;
    8'h2f: p21 <= 8'h15;
    8'h30: p21 <= 8'h04;
    8'h31: p21 <= 8'hc7;
    8'h32: p21 <= 8'h23;
    8'h33: p21 <= 8'hc3;
    8'h34: p21 <= 8'h18;
    8'h35: p21 <= 8'h96;
    8'h36: p21 <= 8'h05;
    8'h37: p21 <= 8'h9a;
    8'h38: p21 <= 8'h07;
    8'h39: p21 <= 8'h12;
    8'h3a: p21 <= 8'h80;
    8'h3b: p21 <= 8'he2;
    8'h3c: p21 <= 8'heb;
    8'h3d: p21 <= 8'h27;
    8'h3e: p21 <= 8'hb2;
    8'h3f: p21 <= 8'h75;
    8'h40: p21 <= 8'h09;
    8'h41: p21 <= 8'h83;
    8'h42: p21 <= 8'h2c;
    8'h43: p21 <= 8'h1a;
    8'h44: p21 <= 8'h1b;
    8'h45: p21 <= 8'h6e;
    8'h46: p21 <= 8'h5a;
    8'h47: p21 <= 8'ha0;
    8'h48: p21 <= 8'h52;
    8'h49: p21 <= 8'h3b;
    8'h4a: p21 <= 8'hd6;
    8'h4b: p21 <= 8'hb3;
    8'h4c: p21 <= 8'h29;
    8'h4d: p21 <= 8'he3;
    8'h4e: p21 <= 8'h2f;
    8'h4f: p21 <= 8'h84;
    8'h50: p21 <= 8'h53;
    8'h51: p21 <= 8'hd1;
    8'h52: p21 <= 8'h00;
    8'h53: p21 <= 8'hed;
    8'h54: p21 <= 8'h20;
    8'h55: p21 <= 8'hfc;
    8'h56: p21 <= 8'hb1;
    8'h57: p21 <= 8'h5b;
    8'h58: p21 <= 8'h6a;
    8'h59: p21 <= 8'hcb;
    8'h5a: p21 <= 8'hbe;
    8'h5b: p21 <= 8'h39;
    8'h5c: p21 <= 8'h4a;
    8'h5d: p21 <= 8'h4c;
    8'h5e: p21 <= 8'h58;
    8'h5f: p21 <= 8'hcf;
    8'h60: p21 <= 8'hd0;
    8'h61: p21 <= 8'hef;
    8'h62: p21 <= 8'haa;
    8'h63: p21 <= 8'hfb;
    8'h64: p21 <= 8'h43;
    8'h65: p21 <= 8'h4d;
    8'h66: p21 <= 8'h33;
    8'h67: p21 <= 8'h85;
    8'h68: p21 <= 8'h45;
    8'h69: p21 <= 8'hf9;
    8'h6a: p21 <= 8'h02;
    8'h6b: p21 <= 8'h7f;
    8'h6c: p21 <= 8'h50;
    8'h6d: p21 <= 8'h3c;
    8'h6e: p21 <= 8'h9f;
    8'h6f: p21 <= 8'ha8;
    8'h70: p21 <= 8'h51;
    8'h71: p21 <= 8'ha3;
    8'h72: p21 <= 8'h40;
    8'h73: p21 <= 8'h8f;
    8'h74: p21 <= 8'h92;
    8'h75: p21 <= 8'h9d;
    8'h76: p21 <= 8'h38;
    8'h77: p21 <= 8'hf5;
    8'h78: p21 <= 8'hbc;
    8'h79: p21 <= 8'hb6;
    8'h7a: p21 <= 8'hda;
    8'h7b: p21 <= 8'h21;
    8'h7c: p21 <= 8'h10;
    8'h7d: p21 <= 8'hff;
    8'h7e: p21 <= 8'hf3;
    8'h7f: p21 <= 8'hd2;
    8'h80: p21 <= 8'hcd;
    8'h81: p21 <= 8'h0c;
    8'h82: p21 <= 8'h13;
    8'h83: p21 <= 8'hec;
    8'h84: p21 <= 8'h5f;
    8'h85: p21 <= 8'h97;
    8'h86: p21 <= 8'h44;
    8'h87: p21 <= 8'h17;
    8'h88: p21 <= 8'hc4;
    8'h89: p21 <= 8'ha7;
    8'h8a: p21 <= 8'h7e;
    8'h8b: p21 <= 8'h3d;
    8'h8c: p21 <= 8'h64;
    8'h8d: p21 <= 8'h5d;
    8'h8e: p21 <= 8'h19;
    8'h8f: p21 <= 8'h73;
    8'h90: p21 <= 8'h60;
    8'h91: p21 <= 8'h81;
    8'h92: p21 <= 8'h4f;
    8'h93: p21 <= 8'hdc;
    8'h94: p21 <= 8'h22;
    8'h95: p21 <= 8'h2a;
    8'h96: p21 <= 8'h90;
    8'h97: p21 <= 8'h88;
    8'h98: p21 <= 8'h46;
    8'h99: p21 <= 8'hee;
    8'h9a: p21 <= 8'hb8;
    8'h9b: p21 <= 8'h14;
    8'h9c: p21 <= 8'hde;
    8'h9d: p21 <= 8'h5e;
    8'h9e: p21 <= 8'h0b;
    8'h9f: p21 <= 8'hdb;
    8'ha0: p21 <= 8'he0;
    8'ha1: p21 <= 8'h32;
    8'ha2: p21 <= 8'h3a;
    8'ha3: p21 <= 8'h0a;
    8'ha4: p21 <= 8'h49;
    8'ha5: p21 <= 8'h06;
    8'ha6: p21 <= 8'h24;
    8'ha7: p21 <= 8'h5c;
    8'ha8: p21 <= 8'hc2;
    8'ha9: p21 <= 8'hd3;
    8'haa: p21 <= 8'hac;
    8'hab: p21 <= 8'h62;
    8'hac: p21 <= 8'h91;
    8'had: p21 <= 8'h95;
    8'hae: p21 <= 8'he4;
    8'haf: p21 <= 8'h79;
    8'hb0: p21 <= 8'he7;
    8'hb1: p21 <= 8'hc8;
    8'hb2: p21 <= 8'h37;
    8'hb3: p21 <= 8'h6d;
    8'hb4: p21 <= 8'h8d;
    8'hb5: p21 <= 8'hd5;
    8'hb6: p21 <= 8'h4e;
    8'hb7: p21 <= 8'ha9;
    8'hb8: p21 <= 8'h6c;
    8'hb9: p21 <= 8'h56;
    8'hba: p21 <= 8'hf4;
    8'hbb: p21 <= 8'hea;
    8'hbc: p21 <= 8'h65;
    8'hbd: p21 <= 8'h7a;
    8'hbe: p21 <= 8'hae;
    8'hbf: p21 <= 8'h08;
    8'hc0: p21 <= 8'hba;
    8'hc1: p21 <= 8'h78;
    8'hc2: p21 <= 8'h25;
    8'hc3: p21 <= 8'h2e;
    8'hc4: p21 <= 8'h1c;
    8'hc5: p21 <= 8'ha6;
    8'hc6: p21 <= 8'hb4;
    8'hc7: p21 <= 8'hc6;
    8'hc8: p21 <= 8'he8;
    8'hc9: p21 <= 8'hdd;
    8'hca: p21 <= 8'h74;
    8'hcb: p21 <= 8'h1f;
    8'hcc: p21 <= 8'h4b;
    8'hcd: p21 <= 8'hbd;
    8'hce: p21 <= 8'h8b;
    8'hcf: p21 <= 8'h8a;
    8'hd0: p21 <= 8'h70;
    8'hd1: p21 <= 8'h3e;
    8'hd2: p21 <= 8'hb5;
    8'hd3: p21 <= 8'h66;
    8'hd4: p21 <= 8'h48;
    8'hd5: p21 <= 8'h03;
    8'hd6: p21 <= 8'hf6;
    8'hd7: p21 <= 8'h0e;
    8'hd8: p21 <= 8'h61;
    8'hd9: p21 <= 8'h35;
    8'hda: p21 <= 8'h57;
    8'hdb: p21 <= 8'hb9;
    8'hdc: p21 <= 8'h86;
    8'hdd: p21 <= 8'hc1;
    8'hde: p21 <= 8'h1d;
    8'hdf: p21 <= 8'h9e;
    8'he0: p21 <= 8'he1;
    8'he1: p21 <= 8'hf8;
    8'he2: p21 <= 8'h98;
    8'he3: p21 <= 8'h11;
    8'he4: p21 <= 8'h69;
    8'he5: p21 <= 8'hd9;
    8'he6: p21 <= 8'h8e;
    8'he7: p21 <= 8'h94;
    8'he8: p21 <= 8'h9b;
    8'he9: p21 <= 8'h1e;
    8'hea: p21 <= 8'h87;
    8'heb: p21 <= 8'he9;
    8'hec: p21 <= 8'hce;
    8'hed: p21 <= 8'h55;
    8'hee: p21 <= 8'h28;
    8'hef: p21 <= 8'hdf;
    8'hf0: p21 <= 8'h8c;
    8'hf1: p21 <= 8'ha1;
    8'hf2: p21 <= 8'h89;
    8'hf3: p21 <= 8'h0d;
    8'hf4: p21 <= 8'hbf;
    8'hf5: p21 <= 8'he6;
    8'hf6: p21 <= 8'h42;
    8'hf7: p21 <= 8'h68;
    8'hf8: p21 <= 8'h41;
    8'hf9: p21 <= 8'h99;
    8'hfa: p21 <= 8'h2d;
    8'hfb: p21 <= 8'h0f;
    8'hfc: p21 <= 8'hb0;
    8'hfd: p21 <= 8'h54;
    8'hfe: p21 <= 8'hbb;
    8'hff: p21 <= 8'h16;
    endcase
	
    // Third Portion
    case (s2[23:16])
    8'h00: p22 <= 8'h63;
    8'h01: p22 <= 8'h7c;
    8'h02: p22 <= 8'h77;
    8'h03: p22 <= 8'h7b;
    8'h04: p22 <= 8'hf2;
    8'h05: p22 <= 8'h6b;
    8'h06: p22 <= 8'h6f;
    8'h07: p22 <= 8'hc5;
    8'h08: p22 <= 8'h30;
    8'h09: p22 <= 8'h01;
    8'h0a: p22 <= 8'h67;
    8'h0b: p22 <= 8'h2b;
    8'h0c: p22 <= 8'hfe;
    8'h0d: p22 <= 8'hd7;
    8'h0e: p22 <= 8'hab;
    8'h0f: p22 <= 8'h76;
    8'h10: p22 <= 8'hca;
    8'h11: p22 <= 8'h82;
    8'h12: p22 <= 8'hc9;
    8'h13: p22 <= 8'h7d;
    8'h14: p22 <= 8'hfa;
    8'h15: p22 <= 8'h59;
    8'h16: p22 <= 8'h47;
    8'h17: p22 <= 8'hf0;
    8'h18: p22 <= 8'had;
    8'h19: p22 <= 8'hd4;
    8'h1a: p22 <= 8'ha2;
    8'h1b: p22 <= 8'haf;
    8'h1c: p22 <= 8'h9c;
    8'h1d: p22 <= 8'ha4;
    8'h1e: p22 <= 8'h72;
    8'h1f: p22 <= 8'hc0;
    8'h20: p22 <= 8'hb7;
    8'h21: p22 <= 8'hfd;
    8'h22: p22 <= 8'h93;
    8'h23: p22 <= 8'h26;
    8'h24: p22 <= 8'h36;
    8'h25: p22 <= 8'h3f;
    8'h26: p22 <= 8'hf7;
    8'h27: p22 <= 8'hcc;
    8'h28: p22 <= 8'h34;
    8'h29: p22 <= 8'ha5;
    8'h2a: p22 <= 8'he5;
    8'h2b: p22 <= 8'hf1;
    8'h2c: p22 <= 8'h71;
    8'h2d: p22 <= 8'hd8;
    8'h2e: p22 <= 8'h31;
    8'h2f: p22 <= 8'h15;
    8'h30: p22 <= 8'h04;
    8'h31: p22 <= 8'hc7;
    8'h32: p22 <= 8'h23;
    8'h33: p22 <= 8'hc3;
    8'h34: p22 <= 8'h18;
    8'h35: p22 <= 8'h96;
    8'h36: p22 <= 8'h05;
    8'h37: p22 <= 8'h9a;
    8'h38: p22 <= 8'h07;
    8'h39: p22 <= 8'h12;
    8'h3a: p22 <= 8'h80;
    8'h3b: p22 <= 8'he2;
    8'h3c: p22 <= 8'heb;
    8'h3d: p22 <= 8'h27;
    8'h3e: p22 <= 8'hb2;
    8'h3f: p22 <= 8'h75;
    8'h40: p22 <= 8'h09;
    8'h41: p22 <= 8'h83;
    8'h42: p22 <= 8'h2c;
    8'h43: p22 <= 8'h1a;
    8'h44: p22 <= 8'h1b;
    8'h45: p22 <= 8'h6e;
    8'h46: p22 <= 8'h5a;
    8'h47: p22 <= 8'ha0;
    8'h48: p22 <= 8'h52;
    8'h49: p22 <= 8'h3b;
    8'h4a: p22 <= 8'hd6;
    8'h4b: p22 <= 8'hb3;
    8'h4c: p22 <= 8'h29;
    8'h4d: p22 <= 8'he3;
    8'h4e: p22 <= 8'h2f;
    8'h4f: p22 <= 8'h84;
    8'h50: p22 <= 8'h53;
    8'h51: p22 <= 8'hd1;
    8'h52: p22 <= 8'h00;
    8'h53: p22 <= 8'hed;
    8'h54: p22 <= 8'h20;
    8'h55: p22 <= 8'hfc;
    8'h56: p22 <= 8'hb1;
    8'h57: p22 <= 8'h5b;
    8'h58: p22 <= 8'h6a;
    8'h59: p22 <= 8'hcb;
    8'h5a: p22 <= 8'hbe;
    8'h5b: p22 <= 8'h39;
    8'h5c: p22 <= 8'h4a;
    8'h5d: p22 <= 8'h4c;
    8'h5e: p22 <= 8'h58;
    8'h5f: p22 <= 8'hcf;
    8'h60: p22 <= 8'hd0;
    8'h61: p22 <= 8'hef;
    8'h62: p22 <= 8'haa;
    8'h63: p22 <= 8'hfb;
    8'h64: p22 <= 8'h43;
    8'h65: p22 <= 8'h4d;
    8'h66: p22 <= 8'h33;
    8'h67: p22 <= 8'h85;
    8'h68: p22 <= 8'h45;
    8'h69: p22 <= 8'hf9;
    8'h6a: p22 <= 8'h02;
    8'h6b: p22 <= 8'h7f;
    8'h6c: p22 <= 8'h50;
    8'h6d: p22 <= 8'h3c;
    8'h6e: p22 <= 8'h9f;
    8'h6f: p22 <= 8'ha8;
    8'h70: p22 <= 8'h51;
    8'h71: p22 <= 8'ha3;
    8'h72: p22 <= 8'h40;
    8'h73: p22 <= 8'h8f;
    8'h74: p22 <= 8'h92;
    8'h75: p22 <= 8'h9d;
    8'h76: p22 <= 8'h38;
    8'h77: p22 <= 8'hf5;
    8'h78: p22 <= 8'hbc;
    8'h79: p22 <= 8'hb6;
    8'h7a: p22 <= 8'hda;
    8'h7b: p22 <= 8'h21;
    8'h7c: p22 <= 8'h10;
    8'h7d: p22 <= 8'hff;
    8'h7e: p22 <= 8'hf3;
    8'h7f: p22 <= 8'hd2;
    8'h80: p22 <= 8'hcd;
    8'h81: p22 <= 8'h0c;
    8'h82: p22 <= 8'h13;
    8'h83: p22 <= 8'hec;
    8'h84: p22 <= 8'h5f;
    8'h85: p22 <= 8'h97;
    8'h86: p22 <= 8'h44;
    8'h87: p22 <= 8'h17;
    8'h88: p22 <= 8'hc4;
    8'h89: p22 <= 8'ha7;
    8'h8a: p22 <= 8'h7e;
    8'h8b: p22 <= 8'h3d;
    8'h8c: p22 <= 8'h64;
    8'h8d: p22 <= 8'h5d;
    8'h8e: p22 <= 8'h19;
    8'h8f: p22 <= 8'h73;
    8'h90: p22 <= 8'h60;
    8'h91: p22 <= 8'h81;
    8'h92: p22 <= 8'h4f;
    8'h93: p22 <= 8'hdc;
    8'h94: p22 <= 8'h22;
    8'h95: p22 <= 8'h2a;
    8'h96: p22 <= 8'h90;
    8'h97: p22 <= 8'h88;
    8'h98: p22 <= 8'h46;
    8'h99: p22 <= 8'hee;
    8'h9a: p22 <= 8'hb8;
    8'h9b: p22 <= 8'h14;
    8'h9c: p22 <= 8'hde;
    8'h9d: p22 <= 8'h5e;
    8'h9e: p22 <= 8'h0b;
    8'h9f: p22 <= 8'hdb;
    8'ha0: p22 <= 8'he0;
    8'ha1: p22 <= 8'h32;
    8'ha2: p22 <= 8'h3a;
    8'ha3: p22 <= 8'h0a;
    8'ha4: p22 <= 8'h49;
    8'ha5: p22 <= 8'h06;
    8'ha6: p22 <= 8'h24;
    8'ha7: p22 <= 8'h5c;
    8'ha8: p22 <= 8'hc2;
    8'ha9: p22 <= 8'hd3;
    8'haa: p22 <= 8'hac;
    8'hab: p22 <= 8'h62;
    8'hac: p22 <= 8'h91;
    8'had: p22 <= 8'h95;
    8'hae: p22 <= 8'he4;
    8'haf: p22 <= 8'h79;
    8'hb0: p22 <= 8'he7;
    8'hb1: p22 <= 8'hc8;
    8'hb2: p22 <= 8'h37;
    8'hb3: p22 <= 8'h6d;
    8'hb4: p22 <= 8'h8d;
    8'hb5: p22 <= 8'hd5;
    8'hb6: p22 <= 8'h4e;
    8'hb7: p22 <= 8'ha9;
    8'hb8: p22 <= 8'h6c;
    8'hb9: p22 <= 8'h56;
    8'hba: p22 <= 8'hf4;
    8'hbb: p22 <= 8'hea;
    8'hbc: p22 <= 8'h65;
    8'hbd: p22 <= 8'h7a;
    8'hbe: p22 <= 8'hae;
    8'hbf: p22 <= 8'h08;
    8'hc0: p22 <= 8'hba;
    8'hc1: p22 <= 8'h78;
    8'hc2: p22 <= 8'h25;
    8'hc3: p22 <= 8'h2e;
    8'hc4: p22 <= 8'h1c;
    8'hc5: p22 <= 8'ha6;
    8'hc6: p22 <= 8'hb4;
    8'hc7: p22 <= 8'hc6;
    8'hc8: p22 <= 8'he8;
    8'hc9: p22 <= 8'hdd;
    8'hca: p22 <= 8'h74;
    8'hcb: p22 <= 8'h1f;
    8'hcc: p22 <= 8'h4b;
    8'hcd: p22 <= 8'hbd;
    8'hce: p22 <= 8'h8b;
    8'hcf: p22 <= 8'h8a;
    8'hd0: p22 <= 8'h70;
    8'hd1: p22 <= 8'h3e;
    8'hd2: p22 <= 8'hb5;
    8'hd3: p22 <= 8'h66;
    8'hd4: p22 <= 8'h48;
    8'hd5: p22 <= 8'h03;
    8'hd6: p22 <= 8'hf6;
    8'hd7: p22 <= 8'h0e;
    8'hd8: p22 <= 8'h61;
    8'hd9: p22 <= 8'h35;
    8'hda: p22 <= 8'h57;
    8'hdb: p22 <= 8'hb9;
    8'hdc: p22 <= 8'h86;
    8'hdd: p22 <= 8'hc1;
    8'hde: p22 <= 8'h1d;
    8'hdf: p22 <= 8'h9e;
    8'he0: p22 <= 8'he1;
    8'he1: p22 <= 8'hf8;
    8'he2: p22 <= 8'h98;
    8'he3: p22 <= 8'h11;
    8'he4: p22 <= 8'h69;
    8'he5: p22 <= 8'hd9;
    8'he6: p22 <= 8'h8e;
    8'he7: p22 <= 8'h94;
    8'he8: p22 <= 8'h9b;
    8'he9: p22 <= 8'h1e;
    8'hea: p22 <= 8'h87;
    8'heb: p22 <= 8'he9;
    8'hec: p22 <= 8'hce;
    8'hed: p22 <= 8'h55;
    8'hee: p22 <= 8'h28;
    8'hef: p22 <= 8'hdf;
    8'hf0: p22 <= 8'h8c;
    8'hf1: p22 <= 8'ha1;
    8'hf2: p22 <= 8'h89;
    8'hf3: p22 <= 8'h0d;
    8'hf4: p22 <= 8'hbf;
    8'hf5: p22 <= 8'he6;
    8'hf6: p22 <= 8'h42;
    8'hf7: p22 <= 8'h68;
    8'hf8: p22 <= 8'h41;
    8'hf9: p22 <= 8'h99;
    8'hfa: p22 <= 8'h2d;
    8'hfb: p22 <= 8'h0f;
    8'hfc: p22 <= 8'hb0;
    8'hfd: p22 <= 8'h54;
    8'hfe: p22 <= 8'hbb;
    8'hff: p22 <= 8'h16;
    endcase
	
    // Fourth Portion
    case (s2[31:24])
    8'h00: p23 <= 8'h63;
    8'h01: p23 <= 8'h7c;
    8'h02: p23 <= 8'h77;
    8'h03: p23 <= 8'h7b;
    8'h04: p23 <= 8'hf2;
    8'h05: p23 <= 8'h6b;
    8'h06: p23 <= 8'h6f;
    8'h07: p23 <= 8'hc5;
    8'h08: p23 <= 8'h30;
    8'h09: p23 <= 8'h01;
    8'h0a: p23 <= 8'h67;
    8'h0b: p23 <= 8'h2b;
    8'h0c: p23 <= 8'hfe;
    8'h0d: p23 <= 8'hd7;
    8'h0e: p23 <= 8'hab;
    8'h0f: p23 <= 8'h76;
    8'h10: p23 <= 8'hca;
    8'h11: p23 <= 8'h82;
    8'h12: p23 <= 8'hc9;
    8'h13: p23 <= 8'h7d;
    8'h14: p23 <= 8'hfa;
    8'h15: p23 <= 8'h59;
    8'h16: p23 <= 8'h47;
    8'h17: p23 <= 8'hf0;
    8'h18: p23 <= 8'had;
    8'h19: p23 <= 8'hd4;
    8'h1a: p23 <= 8'ha2;
    8'h1b: p23 <= 8'haf;
    8'h1c: p23 <= 8'h9c;
    8'h1d: p23 <= 8'ha4;
    8'h1e: p23 <= 8'h72;
    8'h1f: p23 <= 8'hc0;
    8'h20: p23 <= 8'hb7;
    8'h21: p23 <= 8'hfd;
    8'h22: p23 <= 8'h93;
    8'h23: p23 <= 8'h26;
    8'h24: p23 <= 8'h36;
    8'h25: p23 <= 8'h3f;
    8'h26: p23 <= 8'hf7;
    8'h27: p23 <= 8'hcc;
    8'h28: p23 <= 8'h34;
    8'h29: p23 <= 8'ha5;
    8'h2a: p23 <= 8'he5;
    8'h2b: p23 <= 8'hf1;
    8'h2c: p23 <= 8'h71;
    8'h2d: p23 <= 8'hd8;
    8'h2e: p23 <= 8'h31;
    8'h2f: p23 <= 8'h15;
    8'h30: p23 <= 8'h04;
    8'h31: p23 <= 8'hc7;
    8'h32: p23 <= 8'h23;
    8'h33: p23 <= 8'hc3;
    8'h34: p23 <= 8'h18;
    8'h35: p23 <= 8'h96;
    8'h36: p23 <= 8'h05;
    8'h37: p23 <= 8'h9a;
    8'h38: p23 <= 8'h07;
    8'h39: p23 <= 8'h12;
    8'h3a: p23 <= 8'h80;
    8'h3b: p23 <= 8'he2;
    8'h3c: p23 <= 8'heb;
    8'h3d: p23 <= 8'h27;
    8'h3e: p23 <= 8'hb2;
    8'h3f: p23 <= 8'h75;
    8'h40: p23 <= 8'h09;
    8'h41: p23 <= 8'h83;
    8'h42: p23 <= 8'h2c;
    8'h43: p23 <= 8'h1a;
    8'h44: p23 <= 8'h1b;
    8'h45: p23 <= 8'h6e;
    8'h46: p23 <= 8'h5a;
    8'h47: p23 <= 8'ha0;
    8'h48: p23 <= 8'h52;
    8'h49: p23 <= 8'h3b;
    8'h4a: p23 <= 8'hd6;
    8'h4b: p23 <= 8'hb3;
    8'h4c: p23 <= 8'h29;
    8'h4d: p23 <= 8'he3;
    8'h4e: p23 <= 8'h2f;
    8'h4f: p23 <= 8'h84;
    8'h50: p23 <= 8'h53;
    8'h51: p23 <= 8'hd1;
    8'h52: p23 <= 8'h00;
    8'h53: p23 <= 8'hed;
    8'h54: p23 <= 8'h20;
    8'h55: p23 <= 8'hfc;
    8'h56: p23 <= 8'hb1;
    8'h57: p23 <= 8'h5b;
    8'h58: p23 <= 8'h6a;
    8'h59: p23 <= 8'hcb;
    8'h5a: p23 <= 8'hbe;
    8'h5b: p23 <= 8'h39;
    8'h5c: p23 <= 8'h4a;
    8'h5d: p23 <= 8'h4c;
    8'h5e: p23 <= 8'h58;
    8'h5f: p23 <= 8'hcf;
    8'h60: p23 <= 8'hd0;
    8'h61: p23 <= 8'hef;
    8'h62: p23 <= 8'haa;
    8'h63: p23 <= 8'hfb;
    8'h64: p23 <= 8'h43;
    8'h65: p23 <= 8'h4d;
    8'h66: p23 <= 8'h33;
    8'h67: p23 <= 8'h85;
    8'h68: p23 <= 8'h45;
    8'h69: p23 <= 8'hf9;
    8'h6a: p23 <= 8'h02;
    8'h6b: p23 <= 8'h7f;
    8'h6c: p23 <= 8'h50;
    8'h6d: p23 <= 8'h3c;
    8'h6e: p23 <= 8'h9f;
    8'h6f: p23 <= 8'ha8;
    8'h70: p23 <= 8'h51;
    8'h71: p23 <= 8'ha3;
    8'h72: p23 <= 8'h40;
    8'h73: p23 <= 8'h8f;
    8'h74: p23 <= 8'h92;
    8'h75: p23 <= 8'h9d;
    8'h76: p23 <= 8'h38;
    8'h77: p23 <= 8'hf5;
    8'h78: p23 <= 8'hbc;
    8'h79: p23 <= 8'hb6;
    8'h7a: p23 <= 8'hda;
    8'h7b: p23 <= 8'h21;
    8'h7c: p23 <= 8'h10;
    8'h7d: p23 <= 8'hff;
    8'h7e: p23 <= 8'hf3;
    8'h7f: p23 <= 8'hd2;
    8'h80: p23 <= 8'hcd;
    8'h81: p23 <= 8'h0c;
    8'h82: p23 <= 8'h13;
    8'h83: p23 <= 8'hec;
    8'h84: p23 <= 8'h5f;
    8'h85: p23 <= 8'h97;
    8'h86: p23 <= 8'h44;
    8'h87: p23 <= 8'h17;
    8'h88: p23 <= 8'hc4;
    8'h89: p23 <= 8'ha7;
    8'h8a: p23 <= 8'h7e;
    8'h8b: p23 <= 8'h3d;
    8'h8c: p23 <= 8'h64;
    8'h8d: p23 <= 8'h5d;
    8'h8e: p23 <= 8'h19;
    8'h8f: p23 <= 8'h73;
    8'h90: p23 <= 8'h60;
    8'h91: p23 <= 8'h81;
    8'h92: p23 <= 8'h4f;
    8'h93: p23 <= 8'hdc;
    8'h94: p23 <= 8'h22;
    8'h95: p23 <= 8'h2a;
    8'h96: p23 <= 8'h90;
    8'h97: p23 <= 8'h88;
    8'h98: p23 <= 8'h46;
    8'h99: p23 <= 8'hee;
    8'h9a: p23 <= 8'hb8;
    8'h9b: p23 <= 8'h14;
    8'h9c: p23 <= 8'hde;
    8'h9d: p23 <= 8'h5e;
    8'h9e: p23 <= 8'h0b;
    8'h9f: p23 <= 8'hdb;
    8'ha0: p23 <= 8'he0;
    8'ha1: p23 <= 8'h32;
    8'ha2: p23 <= 8'h3a;
    8'ha3: p23 <= 8'h0a;
    8'ha4: p23 <= 8'h49;
    8'ha5: p23 <= 8'h06;
    8'ha6: p23 <= 8'h24;
    8'ha7: p23 <= 8'h5c;
    8'ha8: p23 <= 8'hc2;
    8'ha9: p23 <= 8'hd3;
    8'haa: p23 <= 8'hac;
    8'hab: p23 <= 8'h62;
    8'hac: p23 <= 8'h91;
    8'had: p23 <= 8'h95;
    8'hae: p23 <= 8'he4;
    8'haf: p23 <= 8'h79;
    8'hb0: p23 <= 8'he7;
    8'hb1: p23 <= 8'hc8;
    8'hb2: p23 <= 8'h37;
    8'hb3: p23 <= 8'h6d;
    8'hb4: p23 <= 8'h8d;
    8'hb5: p23 <= 8'hd5;
    8'hb6: p23 <= 8'h4e;
    8'hb7: p23 <= 8'ha9;
    8'hb8: p23 <= 8'h6c;
    8'hb9: p23 <= 8'h56;
    8'hba: p23 <= 8'hf4;
    8'hbb: p23 <= 8'hea;
    8'hbc: p23 <= 8'h65;
    8'hbd: p23 <= 8'h7a;
    8'hbe: p23 <= 8'hae;
    8'hbf: p23 <= 8'h08;
    8'hc0: p23 <= 8'hba;
    8'hc1: p23 <= 8'h78;
    8'hc2: p23 <= 8'h25;
    8'hc3: p23 <= 8'h2e;
    8'hc4: p23 <= 8'h1c;
    8'hc5: p23 <= 8'ha6;
    8'hc6: p23 <= 8'hb4;
    8'hc7: p23 <= 8'hc6;
    8'hc8: p23 <= 8'he8;
    8'hc9: p23 <= 8'hdd;
    8'hca: p23 <= 8'h74;
    8'hcb: p23 <= 8'h1f;
    8'hcc: p23 <= 8'h4b;
    8'hcd: p23 <= 8'hbd;
    8'hce: p23 <= 8'h8b;
    8'hcf: p23 <= 8'h8a;
    8'hd0: p23 <= 8'h70;
    8'hd1: p23 <= 8'h3e;
    8'hd2: p23 <= 8'hb5;
    8'hd3: p23 <= 8'h66;
    8'hd4: p23 <= 8'h48;
    8'hd5: p23 <= 8'h03;
    8'hd6: p23 <= 8'hf6;
    8'hd7: p23 <= 8'h0e;
    8'hd8: p23 <= 8'h61;
    8'hd9: p23 <= 8'h35;
    8'hda: p23 <= 8'h57;
    8'hdb: p23 <= 8'hb9;
    8'hdc: p23 <= 8'h86;
    8'hdd: p23 <= 8'hc1;
    8'hde: p23 <= 8'h1d;
    8'hdf: p23 <= 8'h9e;
    8'he0: p23 <= 8'he1;
    8'he1: p23 <= 8'hf8;
    8'he2: p23 <= 8'h98;
    8'he3: p23 <= 8'h11;
    8'he4: p23 <= 8'h69;
    8'he5: p23 <= 8'hd9;
    8'he6: p23 <= 8'h8e;
    8'he7: p23 <= 8'h94;
    8'he8: p23 <= 8'h9b;
    8'he9: p23 <= 8'h1e;
    8'hea: p23 <= 8'h87;
    8'heb: p23 <= 8'he9;
    8'hec: p23 <= 8'hce;
    8'hed: p23 <= 8'h55;
    8'hee: p23 <= 8'h28;
    8'hef: p23 <= 8'hdf;
    8'hf0: p23 <= 8'h8c;
    8'hf1: p23 <= 8'ha1;
    8'hf2: p23 <= 8'h89;
    8'hf3: p23 <= 8'h0d;
    8'hf4: p23 <= 8'hbf;
    8'hf5: p23 <= 8'he6;
    8'hf6: p23 <= 8'h42;
    8'hf7: p23 <= 8'h68;
    8'hf8: p23 <= 8'h41;
    8'hf9: p23 <= 8'h99;
    8'hfa: p23 <= 8'h2d;
    8'hfb: p23 <= 8'h0f;
    8'hfc: p23 <= 8'hb0;
    8'hfd: p23 <= 8'h54;
    8'hfe: p23 <= 8'hbb;
    8'hff: p23 <= 8'h16;
    endcase
	
	// **************************** PART S3 ****************************
	
    // First Portion
    case (s3[7:0])
    8'h00: p30 <= 8'h63;
    8'h01: p30 <= 8'h7c;
    8'h02: p30 <= 8'h77;
    8'h03: p30 <= 8'h7b;
    8'h04: p30 <= 8'hf2;
    8'h05: p30 <= 8'h6b;
    8'h06: p30 <= 8'h6f;
    8'h07: p30 <= 8'hc5;
    8'h08: p30 <= 8'h30;
    8'h09: p30 <= 8'h01;
    8'h0a: p30 <= 8'h67;
    8'h0b: p30 <= 8'h2b;
    8'h0c: p30 <= 8'hfe;
    8'h0d: p30 <= 8'hd7;
    8'h0e: p30 <= 8'hab;
    8'h0f: p30 <= 8'h76;
    8'h10: p30 <= 8'hca;
    8'h11: p30 <= 8'h82;
    8'h12: p30 <= 8'hc9;
    8'h13: p30 <= 8'h7d;
    8'h14: p30 <= 8'hfa;
    8'h15: p30 <= 8'h59;
    8'h16: p30 <= 8'h47;
    8'h17: p30 <= 8'hf0;
    8'h18: p30 <= 8'had;
    8'h19: p30 <= 8'hd4;
    8'h1a: p30 <= 8'ha2;
    8'h1b: p30 <= 8'haf;
    8'h1c: p30 <= 8'h9c;
    8'h1d: p30 <= 8'ha4;
    8'h1e: p30 <= 8'h72;
    8'h1f: p30 <= 8'hc0;
    8'h20: p30 <= 8'hb7;
    8'h21: p30 <= 8'hfd;
    8'h22: p30 <= 8'h93;
    8'h23: p30 <= 8'h26;
    8'h24: p30 <= 8'h36;
    8'h25: p30 <= 8'h3f;
    8'h26: p30 <= 8'hf7;
    8'h27: p30 <= 8'hcc;
    8'h28: p30 <= 8'h34;
    8'h29: p30 <= 8'ha5;
    8'h2a: p30 <= 8'he5;
    8'h2b: p30 <= 8'hf1;
    8'h2c: p30 <= 8'h71;
    8'h2d: p30 <= 8'hd8;
    8'h2e: p30 <= 8'h31;
    8'h2f: p30 <= 8'h15;
    8'h30: p30 <= 8'h04;
    8'h31: p30 <= 8'hc7;
    8'h32: p30 <= 8'h23;
    8'h33: p30 <= 8'hc3;
    8'h34: p30 <= 8'h18;
    8'h35: p30 <= 8'h96;
    8'h36: p30 <= 8'h05;
    8'h37: p30 <= 8'h9a;
    8'h38: p30 <= 8'h07;
    8'h39: p30 <= 8'h12;
    8'h3a: p30 <= 8'h80;
    8'h3b: p30 <= 8'he2;
    8'h3c: p30 <= 8'heb;
    8'h3d: p30 <= 8'h27;
    8'h3e: p30 <= 8'hb2;
    8'h3f: p30 <= 8'h75;
    8'h40: p30 <= 8'h09;
    8'h41: p30 <= 8'h83;
    8'h42: p30 <= 8'h2c;
    8'h43: p30 <= 8'h1a;
    8'h44: p30 <= 8'h1b;
    8'h45: p30 <= 8'h6e;
    8'h46: p30 <= 8'h5a;
    8'h47: p30 <= 8'ha0;
    8'h48: p30 <= 8'h52;
    8'h49: p30 <= 8'h3b;
    8'h4a: p30 <= 8'hd6;
    8'h4b: p30 <= 8'hb3;
    8'h4c: p30 <= 8'h29;
    8'h4d: p30 <= 8'he3;
    8'h4e: p30 <= 8'h2f;
    8'h4f: p30 <= 8'h84;
    8'h50: p30 <= 8'h53;
    8'h51: p30 <= 8'hd1;
    8'h52: p30 <= 8'h00;
    8'h53: p30 <= 8'hed;
    8'h54: p30 <= 8'h20;
    8'h55: p30 <= 8'hfc;
    8'h56: p30 <= 8'hb1;
    8'h57: p30 <= 8'h5b;
    8'h58: p30 <= 8'h6a;
    8'h59: p30 <= 8'hcb;
    8'h5a: p30 <= 8'hbe;
    8'h5b: p30 <= 8'h39;
    8'h5c: p30 <= 8'h4a;
    8'h5d: p30 <= 8'h4c;
    8'h5e: p30 <= 8'h58;
    8'h5f: p30 <= 8'hcf;
    8'h60: p30 <= 8'hd0;
    8'h61: p30 <= 8'hef;
    8'h62: p30 <= 8'haa;
    8'h63: p30 <= 8'hfb;
    8'h64: p30 <= 8'h43;
    8'h65: p30 <= 8'h4d;
    8'h66: p30 <= 8'h33;
    8'h67: p30 <= 8'h85;
    8'h68: p30 <= 8'h45;
    8'h69: p30 <= 8'hf9;
    8'h6a: p30 <= 8'h02;
    8'h6b: p30 <= 8'h7f;
    8'h6c: p30 <= 8'h50;
    8'h6d: p30 <= 8'h3c;
    8'h6e: p30 <= 8'h9f;
    8'h6f: p30 <= 8'ha8;
    8'h70: p30 <= 8'h51;
    8'h71: p30 <= 8'ha3;
    8'h72: p30 <= 8'h40;
    8'h73: p30 <= 8'h8f;
    8'h74: p30 <= 8'h92;
    8'h75: p30 <= 8'h9d;
    8'h76: p30 <= 8'h38;
    8'h77: p30 <= 8'hf5;
    8'h78: p30 <= 8'hbc;
    8'h79: p30 <= 8'hb6;
    8'h7a: p30 <= 8'hda;
    8'h7b: p30 <= 8'h21;
    8'h7c: p30 <= 8'h10;
    8'h7d: p30 <= 8'hff;
    8'h7e: p30 <= 8'hf3;
    8'h7f: p30 <= 8'hd2;
    8'h80: p30 <= 8'hcd;
    8'h81: p30 <= 8'h0c;
    8'h82: p30 <= 8'h13;
    8'h83: p30 <= 8'hec;
    8'h84: p30 <= 8'h5f;
    8'h85: p30 <= 8'h97;
    8'h86: p30 <= 8'h44;
    8'h87: p30 <= 8'h17;
    8'h88: p30 <= 8'hc4;
    8'h89: p30 <= 8'ha7;
    8'h8a: p30 <= 8'h7e;
    8'h8b: p30 <= 8'h3d;
    8'h8c: p30 <= 8'h64;
    8'h8d: p30 <= 8'h5d;
    8'h8e: p30 <= 8'h19;
    8'h8f: p30 <= 8'h73;
    8'h90: p30 <= 8'h60;
    8'h91: p30 <= 8'h81;
    8'h92: p30 <= 8'h4f;
    8'h93: p30 <= 8'hdc;
    8'h94: p30 <= 8'h22;
    8'h95: p30 <= 8'h2a;
    8'h96: p30 <= 8'h90;
    8'h97: p30 <= 8'h88;
    8'h98: p30 <= 8'h46;
    8'h99: p30 <= 8'hee;
    8'h9a: p30 <= 8'hb8;
    8'h9b: p30 <= 8'h14;
    8'h9c: p30 <= 8'hde;
    8'h9d: p30 <= 8'h5e;
    8'h9e: p30 <= 8'h0b;
    8'h9f: p30 <= 8'hdb;
    8'ha0: p30 <= 8'he0;
    8'ha1: p30 <= 8'h32;
    8'ha2: p30 <= 8'h3a;
    8'ha3: p30 <= 8'h0a;
    8'ha4: p30 <= 8'h49;
    8'ha5: p30 <= 8'h06;
    8'ha6: p30 <= 8'h24;
    8'ha7: p30 <= 8'h5c;
    8'ha8: p30 <= 8'hc2;
    8'ha9: p30 <= 8'hd3;
    8'haa: p30 <= 8'hac;
    8'hab: p30 <= 8'h62;
    8'hac: p30 <= 8'h91;
    8'had: p30 <= 8'h95;
    8'hae: p30 <= 8'he4;
    8'haf: p30 <= 8'h79;
    8'hb0: p30 <= 8'he7;
    8'hb1: p30 <= 8'hc8;
    8'hb2: p30 <= 8'h37;
    8'hb3: p30 <= 8'h6d;
    8'hb4: p30 <= 8'h8d;
    8'hb5: p30 <= 8'hd5;
    8'hb6: p30 <= 8'h4e;
    8'hb7: p30 <= 8'ha9;
    8'hb8: p30 <= 8'h6c;
    8'hb9: p30 <= 8'h56;
    8'hba: p30 <= 8'hf4;
    8'hbb: p30 <= 8'hea;
    8'hbc: p30 <= 8'h65;
    8'hbd: p30 <= 8'h7a;
    8'hbe: p30 <= 8'hae;
    8'hbf: p30 <= 8'h08;
    8'hc0: p30 <= 8'hba;
    8'hc1: p30 <= 8'h78;
    8'hc2: p30 <= 8'h25;
    8'hc3: p30 <= 8'h2e;
    8'hc4: p30 <= 8'h1c;
    8'hc5: p30 <= 8'ha6;
    8'hc6: p30 <= 8'hb4;
    8'hc7: p30 <= 8'hc6;
    8'hc8: p30 <= 8'he8;
    8'hc9: p30 <= 8'hdd;
    8'hca: p30 <= 8'h74;
    8'hcb: p30 <= 8'h1f;
    8'hcc: p30 <= 8'h4b;
    8'hcd: p30 <= 8'hbd;
    8'hce: p30 <= 8'h8b;
    8'hcf: p30 <= 8'h8a;
    8'hd0: p30 <= 8'h70;
    8'hd1: p30 <= 8'h3e;
    8'hd2: p30 <= 8'hb5;
    8'hd3: p30 <= 8'h66;
    8'hd4: p30 <= 8'h48;
    8'hd5: p30 <= 8'h03;
    8'hd6: p30 <= 8'hf6;
    8'hd7: p30 <= 8'h0e;
    8'hd8: p30 <= 8'h61;
    8'hd9: p30 <= 8'h35;
    8'hda: p30 <= 8'h57;
    8'hdb: p30 <= 8'hb9;
    8'hdc: p30 <= 8'h86;
    8'hdd: p30 <= 8'hc1;
    8'hde: p30 <= 8'h1d;
    8'hdf: p30 <= 8'h9e;
    8'he0: p30 <= 8'he1;
    8'he1: p30 <= 8'hf8;
    8'he2: p30 <= 8'h98;
    8'he3: p30 <= 8'h11;
    8'he4: p30 <= 8'h69;
    8'he5: p30 <= 8'hd9;
    8'he6: p30 <= 8'h8e;
    8'he7: p30 <= 8'h94;
    8'he8: p30 <= 8'h9b;
    8'he9: p30 <= 8'h1e;
    8'hea: p30 <= 8'h87;
    8'heb: p30 <= 8'he9;
    8'hec: p30 <= 8'hce;
    8'hed: p30 <= 8'h55;
    8'hee: p30 <= 8'h28;
    8'hef: p30 <= 8'hdf;
    8'hf0: p30 <= 8'h8c;
    8'hf1: p30 <= 8'ha1;
    8'hf2: p30 <= 8'h89;
    8'hf3: p30 <= 8'h0d;
    8'hf4: p30 <= 8'hbf;
    8'hf5: p30 <= 8'he6;
    8'hf6: p30 <= 8'h42;
    8'hf7: p30 <= 8'h68;
    8'hf8: p30 <= 8'h41;
    8'hf9: p30 <= 8'h99;
    8'hfa: p30 <= 8'h2d;
    8'hfb: p30 <= 8'h0f;
    8'hfc: p30 <= 8'hb0;
    8'hfd: p30 <= 8'h54;
    8'hfe: p30 <= 8'hbb;
    8'hff: p30 <= 8'h16;
    endcase
	
    // Second Portion
    case (s3[15:8])
    8'h00: p31 <= 8'h63;
    8'h01: p31 <= 8'h7c;
    8'h02: p31 <= 8'h77;
    8'h03: p31 <= 8'h7b;
    8'h04: p31 <= 8'hf2;
    8'h05: p31 <= 8'h6b;
    8'h06: p31 <= 8'h6f;
    8'h07: p31 <= 8'hc5;
    8'h08: p31 <= 8'h30;
    8'h09: p31 <= 8'h01;
    8'h0a: p31 <= 8'h67;
    8'h0b: p31 <= 8'h2b;
    8'h0c: p31 <= 8'hfe;
    8'h0d: p31 <= 8'hd7;
    8'h0e: p31 <= 8'hab;
    8'h0f: p31 <= 8'h76;
    8'h10: p31 <= 8'hca;
    8'h11: p31 <= 8'h82;
    8'h12: p31 <= 8'hc9;
    8'h13: p31 <= 8'h7d;
    8'h14: p31 <= 8'hfa;
    8'h15: p31 <= 8'h59;
    8'h16: p31 <= 8'h47;
    8'h17: p31 <= 8'hf0;
    8'h18: p31 <= 8'had;
    8'h19: p31 <= 8'hd4;
    8'h1a: p31 <= 8'ha2;
    8'h1b: p31 <= 8'haf;
    8'h1c: p31 <= 8'h9c;
    8'h1d: p31 <= 8'ha4;
    8'h1e: p31 <= 8'h72;
    8'h1f: p31 <= 8'hc0;
    8'h20: p31 <= 8'hb7;
    8'h21: p31 <= 8'hfd;
    8'h22: p31 <= 8'h93;
    8'h23: p31 <= 8'h26;
    8'h24: p31 <= 8'h36;
    8'h25: p31 <= 8'h3f;
    8'h26: p31 <= 8'hf7;
    8'h27: p31 <= 8'hcc;
    8'h28: p31 <= 8'h34;
    8'h29: p31 <= 8'ha5;
    8'h2a: p31 <= 8'he5;
    8'h2b: p31 <= 8'hf1;
    8'h2c: p31 <= 8'h71;
    8'h2d: p31 <= 8'hd8;
    8'h2e: p31 <= 8'h31;
    8'h2f: p31 <= 8'h15;
    8'h30: p31 <= 8'h04;
    8'h31: p31 <= 8'hc7;
    8'h32: p31 <= 8'h23;
    8'h33: p31 <= 8'hc3;
    8'h34: p31 <= 8'h18;
    8'h35: p31 <= 8'h96;
    8'h36: p31 <= 8'h05;
    8'h37: p31 <= 8'h9a;
    8'h38: p31 <= 8'h07;
    8'h39: p31 <= 8'h12;
    8'h3a: p31 <= 8'h80;
    8'h3b: p31 <= 8'he2;
    8'h3c: p31 <= 8'heb;
    8'h3d: p31 <= 8'h27;
    8'h3e: p31 <= 8'hb2;
    8'h3f: p31 <= 8'h75;
    8'h40: p31 <= 8'h09;
    8'h41: p31 <= 8'h83;
    8'h42: p31 <= 8'h2c;
    8'h43: p31 <= 8'h1a;
    8'h44: p31 <= 8'h1b;
    8'h45: p31 <= 8'h6e;
    8'h46: p31 <= 8'h5a;
    8'h47: p31 <= 8'ha0;
    8'h48: p31 <= 8'h52;
    8'h49: p31 <= 8'h3b;
    8'h4a: p31 <= 8'hd6;
    8'h4b: p31 <= 8'hb3;
    8'h4c: p31 <= 8'h29;
    8'h4d: p31 <= 8'he3;
    8'h4e: p31 <= 8'h2f;
    8'h4f: p31 <= 8'h84;
    8'h50: p31 <= 8'h53;
    8'h51: p31 <= 8'hd1;
    8'h52: p31 <= 8'h00;
    8'h53: p31 <= 8'hed;
    8'h54: p31 <= 8'h20;
    8'h55: p31 <= 8'hfc;
    8'h56: p31 <= 8'hb1;
    8'h57: p31 <= 8'h5b;
    8'h58: p31 <= 8'h6a;
    8'h59: p31 <= 8'hcb;
    8'h5a: p31 <= 8'hbe;
    8'h5b: p31 <= 8'h39;
    8'h5c: p31 <= 8'h4a;
    8'h5d: p31 <= 8'h4c;
    8'h5e: p31 <= 8'h58;
    8'h5f: p31 <= 8'hcf;
    8'h60: p31 <= 8'hd0;
    8'h61: p31 <= 8'hef;
    8'h62: p31 <= 8'haa;
    8'h63: p31 <= 8'hfb;
    8'h64: p31 <= 8'h43;
    8'h65: p31 <= 8'h4d;
    8'h66: p31 <= 8'h33;
    8'h67: p31 <= 8'h85;
    8'h68: p31 <= 8'h45;
    8'h69: p31 <= 8'hf9;
    8'h6a: p31 <= 8'h02;
    8'h6b: p31 <= 8'h7f;
    8'h6c: p31 <= 8'h50;
    8'h6d: p31 <= 8'h3c;
    8'h6e: p31 <= 8'h9f;
    8'h6f: p31 <= 8'ha8;
    8'h70: p31 <= 8'h51;
    8'h71: p31 <= 8'ha3;
    8'h72: p31 <= 8'h40;
    8'h73: p31 <= 8'h8f;
    8'h74: p31 <= 8'h92;
    8'h75: p31 <= 8'h9d;
    8'h76: p31 <= 8'h38;
    8'h77: p31 <= 8'hf5;
    8'h78: p31 <= 8'hbc;
    8'h79: p31 <= 8'hb6;
    8'h7a: p31 <= 8'hda;
    8'h7b: p31 <= 8'h21;
    8'h7c: p31 <= 8'h10;
    8'h7d: p31 <= 8'hff;
    8'h7e: p31 <= 8'hf3;
    8'h7f: p31 <= 8'hd2;
    8'h80: p31 <= 8'hcd;
    8'h81: p31 <= 8'h0c;
    8'h82: p31 <= 8'h13;
    8'h83: p31 <= 8'hec;
    8'h84: p31 <= 8'h5f;
    8'h85: p31 <= 8'h97;
    8'h86: p31 <= 8'h44;
    8'h87: p31 <= 8'h17;
    8'h88: p31 <= 8'hc4;
    8'h89: p31 <= 8'ha7;
    8'h8a: p31 <= 8'h7e;
    8'h8b: p31 <= 8'h3d;
    8'h8c: p31 <= 8'h64;
    8'h8d: p31 <= 8'h5d;
    8'h8e: p31 <= 8'h19;
    8'h8f: p31 <= 8'h73;
    8'h90: p31 <= 8'h60;
    8'h91: p31 <= 8'h81;
    8'h92: p31 <= 8'h4f;
    8'h93: p31 <= 8'hdc;
    8'h94: p31 <= 8'h22;
    8'h95: p31 <= 8'h2a;
    8'h96: p31 <= 8'h90;
    8'h97: p31 <= 8'h88;
    8'h98: p31 <= 8'h46;
    8'h99: p31 <= 8'hee;
    8'h9a: p31 <= 8'hb8;
    8'h9b: p31 <= 8'h14;
    8'h9c: p31 <= 8'hde;
    8'h9d: p31 <= 8'h5e;
    8'h9e: p31 <= 8'h0b;
    8'h9f: p31 <= 8'hdb;
    8'ha0: p31 <= 8'he0;
    8'ha1: p31 <= 8'h32;
    8'ha2: p31 <= 8'h3a;
    8'ha3: p31 <= 8'h0a;
    8'ha4: p31 <= 8'h49;
    8'ha5: p31 <= 8'h06;
    8'ha6: p31 <= 8'h24;
    8'ha7: p31 <= 8'h5c;
    8'ha8: p31 <= 8'hc2;
    8'ha9: p31 <= 8'hd3;
    8'haa: p31 <= 8'hac;
    8'hab: p31 <= 8'h62;
    8'hac: p31 <= 8'h91;
    8'had: p31 <= 8'h95;
    8'hae: p31 <= 8'he4;
    8'haf: p31 <= 8'h79;
    8'hb0: p31 <= 8'he7;
    8'hb1: p31 <= 8'hc8;
    8'hb2: p31 <= 8'h37;
    8'hb3: p31 <= 8'h6d;
    8'hb4: p31 <= 8'h8d;
    8'hb5: p31 <= 8'hd5;
    8'hb6: p31 <= 8'h4e;
    8'hb7: p31 <= 8'ha9;
    8'hb8: p31 <= 8'h6c;
    8'hb9: p31 <= 8'h56;
    8'hba: p31 <= 8'hf4;
    8'hbb: p31 <= 8'hea;
    8'hbc: p31 <= 8'h65;
    8'hbd: p31 <= 8'h7a;
    8'hbe: p31 <= 8'hae;
    8'hbf: p31 <= 8'h08;
    8'hc0: p31 <= 8'hba;
    8'hc1: p31 <= 8'h78;
    8'hc2: p31 <= 8'h25;
    8'hc3: p31 <= 8'h2e;
    8'hc4: p31 <= 8'h1c;
    8'hc5: p31 <= 8'ha6;
    8'hc6: p31 <= 8'hb4;
    8'hc7: p31 <= 8'hc6;
    8'hc8: p31 <= 8'he8;
    8'hc9: p31 <= 8'hdd;
    8'hca: p31 <= 8'h74;
    8'hcb: p31 <= 8'h1f;
    8'hcc: p31 <= 8'h4b;
    8'hcd: p31 <= 8'hbd;
    8'hce: p31 <= 8'h8b;
    8'hcf: p31 <= 8'h8a;
    8'hd0: p31 <= 8'h70;
    8'hd1: p31 <= 8'h3e;
    8'hd2: p31 <= 8'hb5;
    8'hd3: p31 <= 8'h66;
    8'hd4: p31 <= 8'h48;
    8'hd5: p31 <= 8'h03;
    8'hd6: p31 <= 8'hf6;
    8'hd7: p31 <= 8'h0e;
    8'hd8: p31 <= 8'h61;
    8'hd9: p31 <= 8'h35;
    8'hda: p31 <= 8'h57;
    8'hdb: p31 <= 8'hb9;
    8'hdc: p31 <= 8'h86;
    8'hdd: p31 <= 8'hc1;
    8'hde: p31 <= 8'h1d;
    8'hdf: p31 <= 8'h9e;
    8'he0: p31 <= 8'he1;
    8'he1: p31 <= 8'hf8;
    8'he2: p31 <= 8'h98;
    8'he3: p31 <= 8'h11;
    8'he4: p31 <= 8'h69;
    8'he5: p31 <= 8'hd9;
    8'he6: p31 <= 8'h8e;
    8'he7: p31 <= 8'h94;
    8'he8: p31 <= 8'h9b;
    8'he9: p31 <= 8'h1e;
    8'hea: p31 <= 8'h87;
    8'heb: p31 <= 8'he9;
    8'hec: p31 <= 8'hce;
    8'hed: p31 <= 8'h55;
    8'hee: p31 <= 8'h28;
    8'hef: p31 <= 8'hdf;
    8'hf0: p31 <= 8'h8c;
    8'hf1: p31 <= 8'ha1;
    8'hf2: p31 <= 8'h89;
    8'hf3: p31 <= 8'h0d;
    8'hf4: p31 <= 8'hbf;
    8'hf5: p31 <= 8'he6;
    8'hf6: p31 <= 8'h42;
    8'hf7: p31 <= 8'h68;
    8'hf8: p31 <= 8'h41;
    8'hf9: p31 <= 8'h99;
    8'hfa: p31 <= 8'h2d;
    8'hfb: p31 <= 8'h0f;
    8'hfc: p31 <= 8'hb0;
    8'hfd: p31 <= 8'h54;
    8'hfe: p31 <= 8'hbb;
    8'hff: p31 <= 8'h16;
    endcase
	
    // Third Portion
    case (s3[23:16])
    8'h00: p32 <= 8'h63;
    8'h01: p32 <= 8'h7c;
    8'h02: p32 <= 8'h77;
    8'h03: p32 <= 8'h7b;
    8'h04: p32 <= 8'hf2;
    8'h05: p32 <= 8'h6b;
    8'h06: p32 <= 8'h6f;
    8'h07: p32 <= 8'hc5;
    8'h08: p32 <= 8'h30;
    8'h09: p32 <= 8'h01;
    8'h0a: p32 <= 8'h67;
    8'h0b: p32 <= 8'h2b;
    8'h0c: p32 <= 8'hfe;
    8'h0d: p32 <= 8'hd7;
    8'h0e: p32 <= 8'hab;
    8'h0f: p32 <= 8'h76;
    8'h10: p32 <= 8'hca;
    8'h11: p32 <= 8'h82;
    8'h12: p32 <= 8'hc9;
    8'h13: p32 <= 8'h7d;
    8'h14: p32 <= 8'hfa;
    8'h15: p32 <= 8'h59;
    8'h16: p32 <= 8'h47;
    8'h17: p32 <= 8'hf0;
    8'h18: p32 <= 8'had;
    8'h19: p32 <= 8'hd4;
    8'h1a: p32 <= 8'ha2;
    8'h1b: p32 <= 8'haf;
    8'h1c: p32 <= 8'h9c;
    8'h1d: p32 <= 8'ha4;
    8'h1e: p32 <= 8'h72;
    8'h1f: p32 <= 8'hc0;
    8'h20: p32 <= 8'hb7;
    8'h21: p32 <= 8'hfd;
    8'h22: p32 <= 8'h93;
    8'h23: p32 <= 8'h26;
    8'h24: p32 <= 8'h36;
    8'h25: p32 <= 8'h3f;
    8'h26: p32 <= 8'hf7;
    8'h27: p32 <= 8'hcc;
    8'h28: p32 <= 8'h34;
    8'h29: p32 <= 8'ha5;
    8'h2a: p32 <= 8'he5;
    8'h2b: p32 <= 8'hf1;
    8'h2c: p32 <= 8'h71;
    8'h2d: p32 <= 8'hd8;
    8'h2e: p32 <= 8'h31;
    8'h2f: p32 <= 8'h15;
    8'h30: p32 <= 8'h04;
    8'h31: p32 <= 8'hc7;
    8'h32: p32 <= 8'h23;
    8'h33: p32 <= 8'hc3;
    8'h34: p32 <= 8'h18;
    8'h35: p32 <= 8'h96;
    8'h36: p32 <= 8'h05;
    8'h37: p32 <= 8'h9a;
    8'h38: p32 <= 8'h07;
    8'h39: p32 <= 8'h12;
    8'h3a: p32 <= 8'h80;
    8'h3b: p32 <= 8'he2;
    8'h3c: p32 <= 8'heb;
    8'h3d: p32 <= 8'h27;
    8'h3e: p32 <= 8'hb2;
    8'h3f: p32 <= 8'h75;
    8'h40: p32 <= 8'h09;
    8'h41: p32 <= 8'h83;
    8'h42: p32 <= 8'h2c;
    8'h43: p32 <= 8'h1a;
    8'h44: p32 <= 8'h1b;
    8'h45: p32 <= 8'h6e;
    8'h46: p32 <= 8'h5a;
    8'h47: p32 <= 8'ha0;
    8'h48: p32 <= 8'h52;
    8'h49: p32 <= 8'h3b;
    8'h4a: p32 <= 8'hd6;
    8'h4b: p32 <= 8'hb3;
    8'h4c: p32 <= 8'h29;
    8'h4d: p32 <= 8'he3;
    8'h4e: p32 <= 8'h2f;
    8'h4f: p32 <= 8'h84;
    8'h50: p32 <= 8'h53;
    8'h51: p32 <= 8'hd1;
    8'h52: p32 <= 8'h00;
    8'h53: p32 <= 8'hed;
    8'h54: p32 <= 8'h20;
    8'h55: p32 <= 8'hfc;
    8'h56: p32 <= 8'hb1;
    8'h57: p32 <= 8'h5b;
    8'h58: p32 <= 8'h6a;
    8'h59: p32 <= 8'hcb;
    8'h5a: p32 <= 8'hbe;
    8'h5b: p32 <= 8'h39;
    8'h5c: p32 <= 8'h4a;
    8'h5d: p32 <= 8'h4c;
    8'h5e: p32 <= 8'h58;
    8'h5f: p32 <= 8'hcf;
    8'h60: p32 <= 8'hd0;
    8'h61: p32 <= 8'hef;
    8'h62: p32 <= 8'haa;
    8'h63: p32 <= 8'hfb;
    8'h64: p32 <= 8'h43;
    8'h65: p32 <= 8'h4d;
    8'h66: p32 <= 8'h33;
    8'h67: p32 <= 8'h85;
    8'h68: p32 <= 8'h45;
    8'h69: p32 <= 8'hf9;
    8'h6a: p32 <= 8'h02;
    8'h6b: p32 <= 8'h7f;
    8'h6c: p32 <= 8'h50;
    8'h6d: p32 <= 8'h3c;
    8'h6e: p32 <= 8'h9f;
    8'h6f: p32 <= 8'ha8;
    8'h70: p32 <= 8'h51;
    8'h71: p32 <= 8'ha3;
    8'h72: p32 <= 8'h40;
    8'h73: p32 <= 8'h8f;
    8'h74: p32 <= 8'h92;
    8'h75: p32 <= 8'h9d;
    8'h76: p32 <= 8'h38;
    8'h77: p32 <= 8'hf5;
    8'h78: p32 <= 8'hbc;
    8'h79: p32 <= 8'hb6;
    8'h7a: p32 <= 8'hda;
    8'h7b: p32 <= 8'h21;
    8'h7c: p32 <= 8'h10;
    8'h7d: p32 <= 8'hff;
    8'h7e: p32 <= 8'hf3;
    8'h7f: p32 <= 8'hd2;
    8'h80: p32 <= 8'hcd;
    8'h81: p32 <= 8'h0c;
    8'h82: p32 <= 8'h13;
    8'h83: p32 <= 8'hec;
    8'h84: p32 <= 8'h5f;
    8'h85: p32 <= 8'h97;
    8'h86: p32 <= 8'h44;
    8'h87: p32 <= 8'h17;
    8'h88: p32 <= 8'hc4;
    8'h89: p32 <= 8'ha7;
    8'h8a: p32 <= 8'h7e;
    8'h8b: p32 <= 8'h3d;
    8'h8c: p32 <= 8'h64;
    8'h8d: p32 <= 8'h5d;
    8'h8e: p32 <= 8'h19;
    8'h8f: p32 <= 8'h73;
    8'h90: p32 <= 8'h60;
    8'h91: p32 <= 8'h81;
    8'h92: p32 <= 8'h4f;
    8'h93: p32 <= 8'hdc;
    8'h94: p32 <= 8'h22;
    8'h95: p32 <= 8'h2a;
    8'h96: p32 <= 8'h90;
    8'h97: p32 <= 8'h88;
    8'h98: p32 <= 8'h46;
    8'h99: p32 <= 8'hee;
    8'h9a: p32 <= 8'hb8;
    8'h9b: p32 <= 8'h14;
    8'h9c: p32 <= 8'hde;
    8'h9d: p32 <= 8'h5e;
    8'h9e: p32 <= 8'h0b;
    8'h9f: p32 <= 8'hdb;
    8'ha0: p32 <= 8'he0;
    8'ha1: p32 <= 8'h32;
    8'ha2: p32 <= 8'h3a;
    8'ha3: p32 <= 8'h0a;
    8'ha4: p32 <= 8'h49;
    8'ha5: p32 <= 8'h06;
    8'ha6: p32 <= 8'h24;
    8'ha7: p32 <= 8'h5c;
    8'ha8: p32 <= 8'hc2;
    8'ha9: p32 <= 8'hd3;
    8'haa: p32 <= 8'hac;
    8'hab: p32 <= 8'h62;
    8'hac: p32 <= 8'h91;
    8'had: p32 <= 8'h95;
    8'hae: p32 <= 8'he4;
    8'haf: p32 <= 8'h79;
    8'hb0: p32 <= 8'he7;
    8'hb1: p32 <= 8'hc8;
    8'hb2: p32 <= 8'h37;
    8'hb3: p32 <= 8'h6d;
    8'hb4: p32 <= 8'h8d;
    8'hb5: p32 <= 8'hd5;
    8'hb6: p32 <= 8'h4e;
    8'hb7: p32 <= 8'ha9;
    8'hb8: p32 <= 8'h6c;
    8'hb9: p32 <= 8'h56;
    8'hba: p32 <= 8'hf4;
    8'hbb: p32 <= 8'hea;
    8'hbc: p32 <= 8'h65;
    8'hbd: p32 <= 8'h7a;
    8'hbe: p32 <= 8'hae;
    8'hbf: p32 <= 8'h08;
    8'hc0: p32 <= 8'hba;
    8'hc1: p32 <= 8'h78;
    8'hc2: p32 <= 8'h25;
    8'hc3: p32 <= 8'h2e;
    8'hc4: p32 <= 8'h1c;
    8'hc5: p32 <= 8'ha6;
    8'hc6: p32 <= 8'hb4;
    8'hc7: p32 <= 8'hc6;
    8'hc8: p32 <= 8'he8;
    8'hc9: p32 <= 8'hdd;
    8'hca: p32 <= 8'h74;
    8'hcb: p32 <= 8'h1f;
    8'hcc: p32 <= 8'h4b;
    8'hcd: p32 <= 8'hbd;
    8'hce: p32 <= 8'h8b;
    8'hcf: p32 <= 8'h8a;
    8'hd0: p32 <= 8'h70;
    8'hd1: p32 <= 8'h3e;
    8'hd2: p32 <= 8'hb5;
    8'hd3: p32 <= 8'h66;
    8'hd4: p32 <= 8'h48;
    8'hd5: p32 <= 8'h03;
    8'hd6: p32 <= 8'hf6;
    8'hd7: p32 <= 8'h0e;
    8'hd8: p32 <= 8'h61;
    8'hd9: p32 <= 8'h35;
    8'hda: p32 <= 8'h57;
    8'hdb: p32 <= 8'hb9;
    8'hdc: p32 <= 8'h86;
    8'hdd: p32 <= 8'hc1;
    8'hde: p32 <= 8'h1d;
    8'hdf: p32 <= 8'h9e;
    8'he0: p32 <= 8'he1;
    8'he1: p32 <= 8'hf8;
    8'he2: p32 <= 8'h98;
    8'he3: p32 <= 8'h11;
    8'he4: p32 <= 8'h69;
    8'he5: p32 <= 8'hd9;
    8'he6: p32 <= 8'h8e;
    8'he7: p32 <= 8'h94;
    8'he8: p32 <= 8'h9b;
    8'he9: p32 <= 8'h1e;
    8'hea: p32 <= 8'h87;
    8'heb: p32 <= 8'he9;
    8'hec: p32 <= 8'hce;
    8'hed: p32 <= 8'h55;
    8'hee: p32 <= 8'h28;
    8'hef: p32 <= 8'hdf;
    8'hf0: p32 <= 8'h8c;
    8'hf1: p32 <= 8'ha1;
    8'hf2: p32 <= 8'h89;
    8'hf3: p32 <= 8'h0d;
    8'hf4: p32 <= 8'hbf;
    8'hf5: p32 <= 8'he6;
    8'hf6: p32 <= 8'h42;
    8'hf7: p32 <= 8'h68;
    8'hf8: p32 <= 8'h41;
    8'hf9: p32 <= 8'h99;
    8'hfa: p32 <= 8'h2d;
    8'hfb: p32 <= 8'h0f;
    8'hfc: p32 <= 8'hb0;
    8'hfd: p32 <= 8'h54;
    8'hfe: p32 <= 8'hbb;
    8'hff: p32 <= 8'h16;
    endcase
	
    // Fourth Portion
    case (s3[31:24])
    8'h00: p33 <= 8'h63;
    8'h01: p33 <= 8'h7c;
    8'h02: p33 <= 8'h77;
    8'h03: p33 <= 8'h7b;
    8'h04: p33 <= 8'hf2;
    8'h05: p33 <= 8'h6b;
    8'h06: p33 <= 8'h6f;
    8'h07: p33 <= 8'hc5;
    8'h08: p33 <= 8'h30;
    8'h09: p33 <= 8'h01;
    8'h0a: p33 <= 8'h67;
    8'h0b: p33 <= 8'h2b;
    8'h0c: p33 <= 8'hfe;
    8'h0d: p33 <= 8'hd7;
    8'h0e: p33 <= 8'hab;
    8'h0f: p33 <= 8'h76;
    8'h10: p33 <= 8'hca;
    8'h11: p33 <= 8'h82;
    8'h12: p33 <= 8'hc9;
    8'h13: p33 <= 8'h7d;
    8'h14: p33 <= 8'hfa;
    8'h15: p33 <= 8'h59;
    8'h16: p33 <= 8'h47;
    8'h17: p33 <= 8'hf0;
    8'h18: p33 <= 8'had;
    8'h19: p33 <= 8'hd4;
    8'h1a: p33 <= 8'ha2;
    8'h1b: p33 <= 8'haf;
    8'h1c: p33 <= 8'h9c;
    8'h1d: p33 <= 8'ha4;
    8'h1e: p33 <= 8'h72;
    8'h1f: p33 <= 8'hc0;
    8'h20: p33 <= 8'hb7;
    8'h21: p33 <= 8'hfd;
    8'h22: p33 <= 8'h93;
    8'h23: p33 <= 8'h26;
    8'h24: p33 <= 8'h36;
    8'h25: p33 <= 8'h3f;
    8'h26: p33 <= 8'hf7;
    8'h27: p33 <= 8'hcc;
    8'h28: p33 <= 8'h34;
    8'h29: p33 <= 8'ha5;
    8'h2a: p33 <= 8'he5;
    8'h2b: p33 <= 8'hf1;
    8'h2c: p33 <= 8'h71;
    8'h2d: p33 <= 8'hd8;
    8'h2e: p33 <= 8'h31;
    8'h2f: p33 <= 8'h15;
    8'h30: p33 <= 8'h04;
    8'h31: p33 <= 8'hc7;
    8'h32: p33 <= 8'h23;
    8'h33: p33 <= 8'hc3;
    8'h34: p33 <= 8'h18;
    8'h35: p33 <= 8'h96;
    8'h36: p33 <= 8'h05;
    8'h37: p33 <= 8'h9a;
    8'h38: p33 <= 8'h07;
    8'h39: p33 <= 8'h12;
    8'h3a: p33 <= 8'h80;
    8'h3b: p33 <= 8'he2;
    8'h3c: p33 <= 8'heb;
    8'h3d: p33 <= 8'h27;
    8'h3e: p33 <= 8'hb2;
    8'h3f: p33 <= 8'h75;
    8'h40: p33 <= 8'h09;
    8'h41: p33 <= 8'h83;
    8'h42: p33 <= 8'h2c;
    8'h43: p33 <= 8'h1a;
    8'h44: p33 <= 8'h1b;
    8'h45: p33 <= 8'h6e;
    8'h46: p33 <= 8'h5a;
    8'h47: p33 <= 8'ha0;
    8'h48: p33 <= 8'h52;
    8'h49: p33 <= 8'h3b;
    8'h4a: p33 <= 8'hd6;
    8'h4b: p33 <= 8'hb3;
    8'h4c: p33 <= 8'h29;
    8'h4d: p33 <= 8'he3;
    8'h4e: p33 <= 8'h2f;
    8'h4f: p33 <= 8'h84;
    8'h50: p33 <= 8'h53;
    8'h51: p33 <= 8'hd1;
    8'h52: p33 <= 8'h00;
    8'h53: p33 <= 8'hed;
    8'h54: p33 <= 8'h20;
    8'h55: p33 <= 8'hfc;
    8'h56: p33 <= 8'hb1;
    8'h57: p33 <= 8'h5b;
    8'h58: p33 <= 8'h6a;
    8'h59: p33 <= 8'hcb;
    8'h5a: p33 <= 8'hbe;
    8'h5b: p33 <= 8'h39;
    8'h5c: p33 <= 8'h4a;
    8'h5d: p33 <= 8'h4c;
    8'h5e: p33 <= 8'h58;
    8'h5f: p33 <= 8'hcf;
    8'h60: p33 <= 8'hd0;
    8'h61: p33 <= 8'hef;
    8'h62: p33 <= 8'haa;
    8'h63: p33 <= 8'hfb;
    8'h64: p33 <= 8'h43;
    8'h65: p33 <= 8'h4d;
    8'h66: p33 <= 8'h33;
    8'h67: p33 <= 8'h85;
    8'h68: p33 <= 8'h45;
    8'h69: p33 <= 8'hf9;
    8'h6a: p33 <= 8'h02;
    8'h6b: p33 <= 8'h7f;
    8'h6c: p33 <= 8'h50;
    8'h6d: p33 <= 8'h3c;
    8'h6e: p33 <= 8'h9f;
    8'h6f: p33 <= 8'ha8;
    8'h70: p33 <= 8'h51;
    8'h71: p33 <= 8'ha3;
    8'h72: p33 <= 8'h40;
    8'h73: p33 <= 8'h8f;
    8'h74: p33 <= 8'h92;
    8'h75: p33 <= 8'h9d;
    8'h76: p33 <= 8'h38;
    8'h77: p33 <= 8'hf5;
    8'h78: p33 <= 8'hbc;
    8'h79: p33 <= 8'hb6;
    8'h7a: p33 <= 8'hda;
    8'h7b: p33 <= 8'h21;
    8'h7c: p33 <= 8'h10;
    8'h7d: p33 <= 8'hff;
    8'h7e: p33 <= 8'hf3;
    8'h7f: p33 <= 8'hd2;
    8'h80: p33 <= 8'hcd;
    8'h81: p33 <= 8'h0c;
    8'h82: p33 <= 8'h13;
    8'h83: p33 <= 8'hec;
    8'h84: p33 <= 8'h5f;
    8'h85: p33 <= 8'h97;
    8'h86: p33 <= 8'h44;
    8'h87: p33 <= 8'h17;
    8'h88: p33 <= 8'hc4;
    8'h89: p33 <= 8'ha7;
    8'h8a: p33 <= 8'h7e;
    8'h8b: p33 <= 8'h3d;
    8'h8c: p33 <= 8'h64;
    8'h8d: p33 <= 8'h5d;
    8'h8e: p33 <= 8'h19;
    8'h8f: p33 <= 8'h73;
    8'h90: p33 <= 8'h60;
    8'h91: p33 <= 8'h81;
    8'h92: p33 <= 8'h4f;
    8'h93: p33 <= 8'hdc;
    8'h94: p33 <= 8'h22;
    8'h95: p33 <= 8'h2a;
    8'h96: p33 <= 8'h90;
    8'h97: p33 <= 8'h88;
    8'h98: p33 <= 8'h46;
    8'h99: p33 <= 8'hee;
    8'h9a: p33 <= 8'hb8;
    8'h9b: p33 <= 8'h14;
    8'h9c: p33 <= 8'hde;
    8'h9d: p33 <= 8'h5e;
    8'h9e: p33 <= 8'h0b;
    8'h9f: p33 <= 8'hdb;
    8'ha0: p33 <= 8'he0;
    8'ha1: p33 <= 8'h32;
    8'ha2: p33 <= 8'h3a;
    8'ha3: p33 <= 8'h0a;
    8'ha4: p33 <= 8'h49;
    8'ha5: p33 <= 8'h06;
    8'ha6: p33 <= 8'h24;
    8'ha7: p33 <= 8'h5c;
    8'ha8: p33 <= 8'hc2;
    8'ha9: p33 <= 8'hd3;
    8'haa: p33 <= 8'hac;
    8'hab: p33 <= 8'h62;
    8'hac: p33 <= 8'h91;
    8'had: p33 <= 8'h95;
    8'hae: p33 <= 8'he4;
    8'haf: p33 <= 8'h79;
    8'hb0: p33 <= 8'he7;
    8'hb1: p33 <= 8'hc8;
    8'hb2: p33 <= 8'h37;
    8'hb3: p33 <= 8'h6d;
    8'hb4: p33 <= 8'h8d;
    8'hb5: p33 <= 8'hd5;
    8'hb6: p33 <= 8'h4e;
    8'hb7: p33 <= 8'ha9;
    8'hb8: p33 <= 8'h6c;
    8'hb9: p33 <= 8'h56;
    8'hba: p33 <= 8'hf4;
    8'hbb: p33 <= 8'hea;
    8'hbc: p33 <= 8'h65;
    8'hbd: p33 <= 8'h7a;
    8'hbe: p33 <= 8'hae;
    8'hbf: p33 <= 8'h08;
    8'hc0: p33 <= 8'hba;
    8'hc1: p33 <= 8'h78;
    8'hc2: p33 <= 8'h25;
    8'hc3: p33 <= 8'h2e;
    8'hc4: p33 <= 8'h1c;
    8'hc5: p33 <= 8'ha6;
    8'hc6: p33 <= 8'hb4;
    8'hc7: p33 <= 8'hc6;
    8'hc8: p33 <= 8'he8;
    8'hc9: p33 <= 8'hdd;
    8'hca: p33 <= 8'h74;
    8'hcb: p33 <= 8'h1f;
    8'hcc: p33 <= 8'h4b;
    8'hcd: p33 <= 8'hbd;
    8'hce: p33 <= 8'h8b;
    8'hcf: p33 <= 8'h8a;
    8'hd0: p33 <= 8'h70;
    8'hd1: p33 <= 8'h3e;
    8'hd2: p33 <= 8'hb5;
    8'hd3: p33 <= 8'h66;
    8'hd4: p33 <= 8'h48;
    8'hd5: p33 <= 8'h03;
    8'hd6: p33 <= 8'hf6;
    8'hd7: p33 <= 8'h0e;
    8'hd8: p33 <= 8'h61;
    8'hd9: p33 <= 8'h35;
    8'hda: p33 <= 8'h57;
    8'hdb: p33 <= 8'hb9;
    8'hdc: p33 <= 8'h86;
    8'hdd: p33 <= 8'hc1;
    8'hde: p33 <= 8'h1d;
    8'hdf: p33 <= 8'h9e;
    8'he0: p33 <= 8'he1;
    8'he1: p33 <= 8'hf8;
    8'he2: p33 <= 8'h98;
    8'he3: p33 <= 8'h11;
    8'he4: p33 <= 8'h69;
    8'he5: p33 <= 8'hd9;
    8'he6: p33 <= 8'h8e;
    8'he7: p33 <= 8'h94;
    8'he8: p33 <= 8'h9b;
    8'he9: p33 <= 8'h1e;
    8'hea: p33 <= 8'h87;
    8'heb: p33 <= 8'he9;
    8'hec: p33 <= 8'hce;
    8'hed: p33 <= 8'h55;
    8'hee: p33 <= 8'h28;
    8'hef: p33 <= 8'hdf;
    8'hf0: p33 <= 8'h8c;
    8'hf1: p33 <= 8'ha1;
    8'hf2: p33 <= 8'h89;
    8'hf3: p33 <= 8'h0d;
    8'hf4: p33 <= 8'hbf;
    8'hf5: p33 <= 8'he6;
    8'hf6: p33 <= 8'h42;
    8'hf7: p33 <= 8'h68;
    8'hf8: p33 <= 8'h41;
    8'hf9: p33 <= 8'h99;
    8'hfa: p33 <= 8'h2d;
    8'hfb: p33 <= 8'h0f;
    8'hfc: p33 <= 8'hb0;
    8'hfd: p33 <= 8'h54;
    8'hfe: p33 <= 8'hbb;
    8'hff: p33 <= 8'h16;
    endcase
	
    end

    assign z0 = {p00, p01, p02, p03} ^ k0;
    assign z1 = {p10, p11, p12, p13} ^ k1;
    assign z2 = {p20, p21, p22, p23} ^ k2;
    assign z3 = {p30, p31, p32, p33} ^ k3;

    assign out = {z0, z1, z2, z3};

endmodule

