
module aes_128 ( clk, state, key, out );
  input [127:0] state;
  input [127:0] key;
  output [127:0] out;
  input clk;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n11, n19, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n31, n39, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n51, n59, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n76, n78, n79, n83, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n96, n104, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n116, n124, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n136, n144, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n156, n164, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n176, n184, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n196, n204, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n216, n224, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n236, n244, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n256, n264, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n276, n284, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n296, n304, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n316, n324, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928;
  wire   [31:0] k3;
  wire   [31:0] k2;
  wire   [31:0] k1;
  wire   [31:0] k0;
  wire   [7:0] p00;
  wire   [7:0] p01;
  wire   [7:0] p02;
  wire   [7:0] p03;
  wire   [7:0] p10;
  wire   [7:0] p11;
  wire   [7:0] p12;
  wire   [7:0] p13;
  wire   [7:0] p20;
  wire   [7:0] p21;
  wire   [7:0] p22;
  wire   [7:0] p23;
  wire   [7:0] p30;
  wire   [7:0] p31;
  wire   [7:0] p32;
  wire   [7:0] p33;

  DFFX1_RVT p32_reg_7_ ( .D(n266), .CLK(clk), .Q(p32[7]) );
  DFFX1_RVT p32_reg_6_ ( .D(n269), .CLK(clk), .Q(p32[6]) );
  DFFX1_RVT p32_reg_5_ ( .D(n270), .CLK(clk), .Q(p32[5]) );
  DFFX1_RVT p32_reg_4_ ( .D(n267), .CLK(clk), .Q(p32[4]) );
  DFFX1_RVT p32_reg_3_ ( .D(n272), .CLK(clk), .Q(p32[3]) );
  DFFX1_RVT p32_reg_2_ ( .D(n268), .CLK(clk), .Q(p32[2]) );
  DFFX1_RVT p32_reg_1_ ( .D(n271), .CLK(clk), .Q(p32[1]) );
  DFFX1_RVT p32_reg_0_ ( .D(n273), .CLK(clk), .Q(p32[0]) );
  DFFX1_RVT k0_reg_31_ ( .D(key[127]), .CLK(clk), .Q(k0[31]) );
  DFFX1_RVT k0_reg_30_ ( .D(key[126]), .CLK(clk), .Q(k0[30]) );
  DFFX1_RVT k0_reg_29_ ( .D(key[125]), .CLK(clk), .Q(k0[29]) );
  DFFX1_RVT k0_reg_28_ ( .D(key[124]), .CLK(clk), .Q(k0[28]) );
  DFFX1_RVT k0_reg_27_ ( .D(key[123]), .CLK(clk), .Q(k0[27]) );
  DFFX1_RVT k0_reg_26_ ( .D(key[122]), .CLK(clk), .Q(k0[26]) );
  DFFX1_RVT k0_reg_25_ ( .D(key[121]), .CLK(clk), .Q(k0[25]) );
  DFFX1_RVT k0_reg_24_ ( .D(key[120]), .CLK(clk), .Q(k0[24]) );
  DFFX1_RVT k0_reg_23_ ( .D(key[119]), .CLK(clk), .Q(k0[23]) );
  DFFX1_RVT k0_reg_22_ ( .D(key[118]), .CLK(clk), .Q(k0[22]) );
  DFFX1_RVT k0_reg_21_ ( .D(key[117]), .CLK(clk), .Q(k0[21]) );
  DFFX1_RVT k0_reg_20_ ( .D(key[116]), .CLK(clk), .Q(k0[20]) );
  DFFX1_RVT k0_reg_19_ ( .D(key[115]), .CLK(clk), .Q(k0[19]) );
  DFFX1_RVT k0_reg_18_ ( .D(key[114]), .CLK(clk), .Q(k0[18]) );
  DFFX1_RVT k0_reg_17_ ( .D(key[113]), .CLK(clk), .Q(k0[17]) );
  DFFX1_RVT k0_reg_16_ ( .D(key[112]), .CLK(clk), .Q(k0[16]) );
  DFFX1_RVT k0_reg_15_ ( .D(key[111]), .CLK(clk), .Q(k0[15]) );
  DFFX1_RVT k0_reg_14_ ( .D(key[110]), .CLK(clk), .Q(k0[14]) );
  DFFX1_RVT k0_reg_13_ ( .D(key[109]), .CLK(clk), .Q(k0[13]) );
  DFFX1_RVT k0_reg_12_ ( .D(key[108]), .CLK(clk), .Q(k0[12]) );
  DFFX1_RVT k0_reg_11_ ( .D(key[107]), .CLK(clk), .Q(k0[11]) );
  DFFX1_RVT k0_reg_10_ ( .D(key[106]), .CLK(clk), .Q(k0[10]) );
  DFFX1_RVT k0_reg_9_ ( .D(key[105]), .CLK(clk), .Q(k0[9]) );
  DFFX1_RVT k0_reg_8_ ( .D(key[104]), .CLK(clk), .Q(k0[8]) );
  DFFX1_RVT k0_reg_7_ ( .D(key[103]), .CLK(clk), .Q(k0[7]) );
  DFFX1_RVT k0_reg_6_ ( .D(key[102]), .CLK(clk), .Q(k0[6]) );
  DFFX1_RVT k0_reg_5_ ( .D(key[101]), .CLK(clk), .Q(k0[5]) );
  DFFX1_RVT k0_reg_4_ ( .D(key[100]), .CLK(clk), .Q(k0[4]) );
  DFFX1_RVT k0_reg_3_ ( .D(key[99]), .CLK(clk), .Q(k0[3]) );
  DFFX1_RVT k0_reg_2_ ( .D(key[98]), .CLK(clk), .Q(k0[2]) );
  DFFX1_RVT k0_reg_1_ ( .D(key[97]), .CLK(clk), .Q(k0[1]) );
  DFFX1_RVT k0_reg_0_ ( .D(key[96]), .CLK(clk), .Q(k0[0]) );
  DFFX1_RVT k3_reg_31_ ( .D(key[31]), .CLK(clk), .Q(k3[31]) );
  DFFX1_RVT k3_reg_30_ ( .D(key[30]), .CLK(clk), .Q(k3[30]) );
  DFFX1_RVT k3_reg_29_ ( .D(key[29]), .CLK(clk), .Q(k3[29]) );
  DFFX1_RVT k3_reg_28_ ( .D(key[28]), .CLK(clk), .Q(k3[28]) );
  DFFX1_RVT k3_reg_27_ ( .D(key[27]), .CLK(clk), .Q(k3[27]) );
  DFFX1_RVT k3_reg_26_ ( .D(key[26]), .CLK(clk), .Q(k3[26]) );
  DFFX1_RVT k3_reg_25_ ( .D(key[25]), .CLK(clk), .Q(k3[25]) );
  DFFX1_RVT k3_reg_24_ ( .D(key[24]), .CLK(clk), .Q(k3[24]) );
  DFFX1_RVT k3_reg_23_ ( .D(key[23]), .CLK(clk), .Q(k3[23]) );
  DFFX1_RVT k3_reg_22_ ( .D(key[22]), .CLK(clk), .Q(k3[22]) );
  DFFX1_RVT k3_reg_21_ ( .D(key[21]), .CLK(clk), .Q(k3[21]) );
  DFFX1_RVT k3_reg_20_ ( .D(key[20]), .CLK(clk), .Q(k3[20]) );
  DFFX1_RVT k3_reg_19_ ( .D(key[19]), .CLK(clk), .Q(k3[19]) );
  DFFX1_RVT k3_reg_18_ ( .D(key[18]), .CLK(clk), .Q(k3[18]) );
  DFFX1_RVT k3_reg_17_ ( .D(key[17]), .CLK(clk), .Q(k3[17]) );
  DFFX1_RVT k3_reg_16_ ( .D(key[16]), .CLK(clk), .Q(k3[16]) );
  DFFX1_RVT k3_reg_15_ ( .D(key[15]), .CLK(clk), .Q(k3[15]) );
  DFFX1_RVT k3_reg_14_ ( .D(key[14]), .CLK(clk), .Q(k3[14]) );
  DFFX1_RVT k3_reg_13_ ( .D(key[13]), .CLK(clk), .Q(k3[13]) );
  DFFX1_RVT k3_reg_12_ ( .D(key[12]), .CLK(clk), .Q(k3[12]) );
  DFFX1_RVT k3_reg_11_ ( .D(key[11]), .CLK(clk), .Q(k3[11]) );
  DFFX1_RVT k3_reg_10_ ( .D(key[10]), .CLK(clk), .Q(k3[10]) );
  DFFX1_RVT k3_reg_9_ ( .D(key[9]), .CLK(clk), .Q(k3[9]) );
  DFFX1_RVT k3_reg_8_ ( .D(key[8]), .CLK(clk), .Q(k3[8]) );
  DFFX1_RVT k3_reg_7_ ( .D(key[7]), .CLK(clk), .Q(k3[7]) );
  DFFX1_RVT k3_reg_6_ ( .D(key[6]), .CLK(clk), .Q(k3[6]) );
  DFFX1_RVT k3_reg_5_ ( .D(key[5]), .CLK(clk), .Q(k3[5]) );
  DFFX1_RVT k3_reg_4_ ( .D(key[4]), .CLK(clk), .Q(k3[4]) );
  DFFX1_RVT k3_reg_3_ ( .D(key[3]), .CLK(clk), .Q(k3[3]) );
  DFFX1_RVT k3_reg_2_ ( .D(key[2]), .CLK(clk), .Q(k3[2]) );
  DFFX1_RVT k3_reg_1_ ( .D(key[1]), .CLK(clk), .Q(k3[1]) );
  DFFX1_RVT k3_reg_0_ ( .D(key[0]), .CLK(clk), .Q(k3[0]) );
  DFFX1_RVT p00_reg_7_ ( .D(n62), .CLK(clk), .Q(p00[7]) );
  DFFX1_RVT p00_reg_6_ ( .D(n61), .CLK(clk), .Q(p00[6]) );
  DFFX1_RVT p00_reg_5_ ( .D(n63), .CLK(clk), .Q(p00[5]) );
  DFFX1_RVT p00_reg_4_ ( .D(n64), .CLK(clk), .Q(p00[4]) );
  DFFX1_RVT p00_reg_3_ ( .D(n68), .CLK(clk), .Q(p00[3]) );
  DFFX1_RVT p00_reg_2_ ( .D(n65), .CLK(clk), .Q(p00[2]) );
  DFFX1_RVT p00_reg_1_ ( .D(n66), .CLK(clk), .Q(p00[1]) );
  DFFX1_RVT p00_reg_0_ ( .D(n67), .CLK(clk), .Q(p00[0]) );
  DFFX1_RVT p12_reg_7_ ( .D(n106), .CLK(clk), .Q(p12[7]) );
  DFFX1_RVT p12_reg_6_ ( .D(n109), .CLK(clk), .Q(p12[6]) );
  DFFX1_RVT p12_reg_5_ ( .D(n110), .CLK(clk), .Q(p12[5]) );
  DFFX1_RVT p12_reg_4_ ( .D(n107), .CLK(clk), .Q(p12[4]) );
  DFFX1_RVT p12_reg_3_ ( .D(n112), .CLK(clk), .Q(p12[3]) );
  DFFX1_RVT p12_reg_2_ ( .D(n108), .CLK(clk), .Q(p12[2]) );
  DFFX1_RVT p12_reg_1_ ( .D(n111), .CLK(clk), .Q(p12[1]) );
  DFFX1_RVT p12_reg_0_ ( .D(n113), .CLK(clk), .Q(p12[0]) );
  DFFX1_RVT p21_reg_7_ ( .D(n206), .CLK(clk), .Q(p21[7]) );
  DFFX1_RVT p21_reg_6_ ( .D(n209), .CLK(clk), .Q(p21[6]) );
  DFFX1_RVT p21_reg_5_ ( .D(n210), .CLK(clk), .Q(p21[5]) );
  DFFX1_RVT p21_reg_4_ ( .D(n207), .CLK(clk), .Q(p21[4]) );
  DFFX1_RVT p21_reg_3_ ( .D(n212), .CLK(clk), .Q(p21[3]) );
  DFFX1_RVT p21_reg_2_ ( .D(n208), .CLK(clk), .Q(p21[2]) );
  DFFX1_RVT p21_reg_1_ ( .D(n211), .CLK(clk), .Q(p21[1]) );
  DFFX1_RVT p21_reg_0_ ( .D(n213), .CLK(clk), .Q(p21[0]) );
  DFFX1_RVT p31_reg_7_ ( .D(n286), .CLK(clk), .Q(p31[7]) );
  DFFX1_RVT p31_reg_6_ ( .D(n289), .CLK(clk), .Q(p31[6]) );
  DFFX1_RVT p31_reg_5_ ( .D(n290), .CLK(clk), .Q(p31[5]) );
  DFFX1_RVT p31_reg_4_ ( .D(n287), .CLK(clk), .Q(p31[4]) );
  DFFX1_RVT p31_reg_3_ ( .D(n292), .CLK(clk), .Q(p31[3]) );
  DFFX1_RVT p31_reg_2_ ( .D(n288), .CLK(clk), .Q(p31[2]) );
  DFFX1_RVT p31_reg_1_ ( .D(n291), .CLK(clk), .Q(p31[1]) );
  DFFX1_RVT p31_reg_0_ ( .D(n293), .CLK(clk), .Q(p31[0]) );
  DFFX1_RVT p02_reg_7_ ( .D(n21), .CLK(clk), .Q(p02[7]) );
  DFFX1_RVT p02_reg_6_ ( .D(n24), .CLK(clk), .Q(p02[6]) );
  DFFX1_RVT p02_reg_5_ ( .D(n25), .CLK(clk), .Q(p02[5]) );
  DFFX1_RVT p02_reg_4_ ( .D(n22), .CLK(clk), .Q(p02[4]) );
  DFFX1_RVT p02_reg_3_ ( .D(n27), .CLK(clk), .Q(p02[3]) );
  DFFX1_RVT p02_reg_2_ ( .D(n23), .CLK(clk), .Q(p02[2]) );
  DFFX1_RVT p02_reg_1_ ( .D(n26), .CLK(clk), .Q(p02[1]) );
  DFFX1_RVT p02_reg_0_ ( .D(n28), .CLK(clk), .Q(p02[0]) );
  DFFX1_RVT p22_reg_7_ ( .D(n186), .CLK(clk), .Q(p22[7]) );
  DFFX1_RVT p22_reg_6_ ( .D(n189), .CLK(clk), .Q(p22[6]) );
  DFFX1_RVT p22_reg_5_ ( .D(n190), .CLK(clk), .Q(p22[5]) );
  DFFX1_RVT p22_reg_4_ ( .D(n187), .CLK(clk), .Q(p22[4]) );
  DFFX1_RVT p22_reg_3_ ( .D(n192), .CLK(clk), .Q(p22[3]) );
  DFFX1_RVT p22_reg_2_ ( .D(n188), .CLK(clk), .Q(p22[2]) );
  DFFX1_RVT p22_reg_1_ ( .D(n191), .CLK(clk), .Q(p22[1]) );
  DFFX1_RVT p22_reg_0_ ( .D(n193), .CLK(clk), .Q(p22[0]) );
  DFFX1_RVT p11_reg_7_ ( .D(n126), .CLK(clk), .Q(p11[7]) );
  DFFX1_RVT p11_reg_6_ ( .D(n129), .CLK(clk), .Q(p11[6]) );
  DFFX1_RVT p11_reg_5_ ( .D(n130), .CLK(clk), .Q(p11[5]) );
  DFFX1_RVT p11_reg_4_ ( .D(n127), .CLK(clk), .Q(p11[4]) );
  DFFX1_RVT p11_reg_3_ ( .D(n132), .CLK(clk), .Q(p11[3]) );
  DFFX1_RVT p11_reg_2_ ( .D(n128), .CLK(clk), .Q(p11[2]) );
  DFFX1_RVT p11_reg_1_ ( .D(n131), .CLK(clk), .Q(p11[1]) );
  DFFX1_RVT p11_reg_0_ ( .D(n133), .CLK(clk), .Q(p11[0]) );
  DFFX1_RVT p23_reg_7_ ( .D(n166), .CLK(clk), .Q(p23[7]) );
  DFFX1_RVT p23_reg_6_ ( .D(n169), .CLK(clk), .Q(p23[6]) );
  DFFX1_RVT p23_reg_5_ ( .D(n170), .CLK(clk), .Q(p23[5]) );
  DFFX1_RVT p23_reg_4_ ( .D(n167), .CLK(clk), .Q(p23[4]) );
  DFFX1_RVT p23_reg_3_ ( .D(n172), .CLK(clk), .Q(p23[3]) );
  DFFX1_RVT p23_reg_2_ ( .D(n168), .CLK(clk), .Q(p23[2]) );
  DFFX1_RVT p23_reg_1_ ( .D(n171), .CLK(clk), .Q(p23[1]) );
  DFFX1_RVT p23_reg_0_ ( .D(n173), .CLK(clk), .Q(p23[0]) );
  DFFX1_RVT p20_reg_7_ ( .D(n226), .CLK(clk), .Q(p20[7]) );
  DFFX1_RVT p20_reg_6_ ( .D(n229), .CLK(clk), .Q(p20[6]) );
  DFFX1_RVT p20_reg_5_ ( .D(n230), .CLK(clk), .Q(p20[5]) );
  DFFX1_RVT p20_reg_4_ ( .D(n227), .CLK(clk), .Q(p20[4]) );
  DFFX1_RVT p20_reg_3_ ( .D(n232), .CLK(clk), .Q(p20[3]) );
  DFFX1_RVT p20_reg_2_ ( .D(n228), .CLK(clk), .Q(p20[2]) );
  DFFX1_RVT p20_reg_1_ ( .D(n231), .CLK(clk), .Q(p20[1]) );
  DFFX1_RVT p20_reg_0_ ( .D(n233), .CLK(clk), .Q(p20[0]) );
  DFFX1_RVT p30_reg_7_ ( .D(n306), .CLK(clk), .Q(p30[7]) );
  DFFX1_RVT p30_reg_6_ ( .D(n309), .CLK(clk), .Q(p30[6]) );
  DFFX1_RVT p30_reg_5_ ( .D(n310), .CLK(clk), .Q(p30[5]) );
  DFFX1_RVT p30_reg_4_ ( .D(n307), .CLK(clk), .Q(p30[4]) );
  DFFX1_RVT p30_reg_3_ ( .D(n312), .CLK(clk), .Q(p30[3]) );
  DFFX1_RVT p30_reg_2_ ( .D(n308), .CLK(clk), .Q(p30[2]) );
  DFFX1_RVT p30_reg_1_ ( .D(n311), .CLK(clk), .Q(p30[1]) );
  DFFX1_RVT p30_reg_0_ ( .D(n313), .CLK(clk), .Q(p30[0]) );
  DFFX1_RVT p01_reg_7_ ( .D(n41), .CLK(clk), .Q(p01[7]) );
  DFFX1_RVT p01_reg_6_ ( .D(n44), .CLK(clk), .Q(p01[6]) );
  DFFX1_RVT p01_reg_5_ ( .D(n45), .CLK(clk), .Q(p01[5]) );
  DFFX1_RVT p01_reg_4_ ( .D(n42), .CLK(clk), .Q(p01[4]) );
  DFFX1_RVT p01_reg_3_ ( .D(n47), .CLK(clk), .Q(p01[3]) );
  DFFX1_RVT p01_reg_2_ ( .D(n43), .CLK(clk), .Q(p01[2]) );
  DFFX1_RVT p01_reg_1_ ( .D(n46), .CLK(clk), .Q(p01[1]) );
  DFFX1_RVT p01_reg_0_ ( .D(n48), .CLK(clk), .Q(p01[0]) );
  DFFX1_RVT p10_reg_7_ ( .D(n146), .CLK(clk), .Q(p10[7]) );
  DFFX1_RVT p10_reg_6_ ( .D(n149), .CLK(clk), .Q(p10[6]) );
  DFFX1_RVT p10_reg_5_ ( .D(n150), .CLK(clk), .Q(p10[5]) );
  DFFX1_RVT p10_reg_4_ ( .D(n147), .CLK(clk), .Q(p10[4]) );
  DFFX1_RVT p10_reg_3_ ( .D(n152), .CLK(clk), .Q(p10[3]) );
  DFFX1_RVT p10_reg_2_ ( .D(n148), .CLK(clk), .Q(p10[2]) );
  DFFX1_RVT p10_reg_1_ ( .D(n151), .CLK(clk), .Q(p10[1]) );
  DFFX1_RVT p10_reg_0_ ( .D(n153), .CLK(clk), .Q(p10[0]) );
  DFFX1_RVT k1_reg_31_ ( .D(key[95]), .CLK(clk), .Q(k1[31]) );
  DFFX1_RVT k1_reg_30_ ( .D(key[94]), .CLK(clk), .Q(k1[30]) );
  DFFX1_RVT k1_reg_29_ ( .D(key[93]), .CLK(clk), .Q(k1[29]) );
  DFFX1_RVT k1_reg_28_ ( .D(key[92]), .CLK(clk), .Q(k1[28]) );
  DFFX1_RVT k1_reg_27_ ( .D(key[91]), .CLK(clk), .Q(k1[27]) );
  DFFX1_RVT k1_reg_26_ ( .D(key[90]), .CLK(clk), .Q(k1[26]) );
  DFFX1_RVT k1_reg_25_ ( .D(key[89]), .CLK(clk), .Q(k1[25]) );
  DFFX1_RVT k1_reg_24_ ( .D(key[88]), .CLK(clk), .Q(k1[24]) );
  DFFX1_RVT k1_reg_23_ ( .D(key[87]), .CLK(clk), .Q(k1[23]) );
  DFFX1_RVT k1_reg_22_ ( .D(key[86]), .CLK(clk), .Q(k1[22]) );
  DFFX1_RVT k1_reg_21_ ( .D(key[85]), .CLK(clk), .Q(k1[21]) );
  DFFX1_RVT k1_reg_20_ ( .D(key[84]), .CLK(clk), .Q(k1[20]) );
  DFFX1_RVT k1_reg_19_ ( .D(key[83]), .CLK(clk), .Q(k1[19]) );
  DFFX1_RVT k1_reg_18_ ( .D(key[82]), .CLK(clk), .Q(k1[18]) );
  DFFX1_RVT k1_reg_17_ ( .D(key[81]), .CLK(clk), .Q(k1[17]) );
  DFFX1_RVT k1_reg_16_ ( .D(key[80]), .CLK(clk), .Q(k1[16]) );
  DFFX1_RVT k1_reg_15_ ( .D(key[79]), .CLK(clk), .Q(k1[15]) );
  DFFX1_RVT k1_reg_14_ ( .D(key[78]), .CLK(clk), .Q(k1[14]) );
  DFFX1_RVT k1_reg_13_ ( .D(key[77]), .CLK(clk), .Q(k1[13]) );
  DFFX1_RVT k1_reg_12_ ( .D(key[76]), .CLK(clk), .Q(k1[12]) );
  DFFX1_RVT k1_reg_11_ ( .D(key[75]), .CLK(clk), .Q(k1[11]) );
  DFFX1_RVT k1_reg_10_ ( .D(key[74]), .CLK(clk), .Q(k1[10]) );
  DFFX1_RVT k1_reg_9_ ( .D(key[73]), .CLK(clk), .Q(k1[9]) );
  DFFX1_RVT k1_reg_8_ ( .D(key[72]), .CLK(clk), .Q(k1[8]) );
  DFFX1_RVT k1_reg_7_ ( .D(key[71]), .CLK(clk), .Q(k1[7]) );
  DFFX1_RVT k1_reg_6_ ( .D(key[70]), .CLK(clk), .Q(k1[6]) );
  DFFX1_RVT k1_reg_5_ ( .D(key[69]), .CLK(clk), .Q(k1[5]) );
  DFFX1_RVT k1_reg_4_ ( .D(key[68]), .CLK(clk), .Q(k1[4]) );
  DFFX1_RVT k1_reg_3_ ( .D(key[67]), .CLK(clk), .Q(k1[3]) );
  DFFX1_RVT k1_reg_2_ ( .D(key[66]), .CLK(clk), .Q(k1[2]) );
  DFFX1_RVT k1_reg_1_ ( .D(key[65]), .CLK(clk), .Q(k1[1]) );
  DFFX1_RVT k1_reg_0_ ( .D(key[64]), .CLK(clk), .Q(k1[0]) );
  DFFX1_RVT p13_reg_7_ ( .D(n86), .CLK(clk), .Q(p13[7]) );
  DFFX1_RVT p13_reg_6_ ( .D(n89), .CLK(clk), .Q(p13[6]) );
  DFFX1_RVT p13_reg_5_ ( .D(n90), .CLK(clk), .Q(p13[5]) );
  DFFX1_RVT p13_reg_4_ ( .D(n87), .CLK(clk), .Q(p13[4]) );
  DFFX1_RVT p13_reg_3_ ( .D(n92), .CLK(clk), .Q(p13[3]) );
  DFFX1_RVT p13_reg_2_ ( .D(n88), .CLK(clk), .Q(p13[2]) );
  DFFX1_RVT p13_reg_1_ ( .D(n91), .CLK(clk), .Q(p13[1]) );
  DFFX1_RVT p13_reg_0_ ( .D(n93), .CLK(clk), .Q(p13[0]) );
  DFFX1_RVT p33_reg_7_ ( .D(n246), .CLK(clk), .Q(p33[7]) );
  DFFX1_RVT p33_reg_6_ ( .D(n249), .CLK(clk), .Q(p33[6]) );
  DFFX1_RVT p33_reg_5_ ( .D(n250), .CLK(clk), .Q(p33[5]) );
  DFFX1_RVT p33_reg_4_ ( .D(n247), .CLK(clk), .Q(p33[4]) );
  DFFX1_RVT p33_reg_3_ ( .D(n252), .CLK(clk), .Q(p33[3]) );
  DFFX1_RVT p33_reg_2_ ( .D(n248), .CLK(clk), .Q(p33[2]) );
  DFFX1_RVT p33_reg_1_ ( .D(n251), .CLK(clk), .Q(p33[1]) );
  DFFX1_RVT p33_reg_0_ ( .D(n253), .CLK(clk), .Q(p33[0]) );
  DFFX1_RVT k2_reg_31_ ( .D(key[63]), .CLK(clk), .Q(k2[31]) );
  DFFX1_RVT k2_reg_30_ ( .D(key[62]), .CLK(clk), .Q(k2[30]) );
  DFFX1_RVT k2_reg_29_ ( .D(key[61]), .CLK(clk), .Q(k2[29]) );
  DFFX1_RVT k2_reg_28_ ( .D(key[60]), .CLK(clk), .Q(k2[28]) );
  DFFX1_RVT k2_reg_27_ ( .D(key[59]), .CLK(clk), .Q(k2[27]) );
  DFFX1_RVT k2_reg_26_ ( .D(key[58]), .CLK(clk), .Q(k2[26]) );
  DFFX1_RVT k2_reg_25_ ( .D(key[57]), .CLK(clk), .Q(k2[25]) );
  DFFX1_RVT k2_reg_24_ ( .D(key[56]), .CLK(clk), .Q(k2[24]) );
  DFFX1_RVT k2_reg_23_ ( .D(key[55]), .CLK(clk), .Q(k2[23]) );
  DFFX1_RVT k2_reg_22_ ( .D(key[54]), .CLK(clk), .Q(k2[22]) );
  DFFX1_RVT k2_reg_21_ ( .D(key[53]), .CLK(clk), .Q(k2[21]) );
  DFFX1_RVT k2_reg_20_ ( .D(key[52]), .CLK(clk), .Q(k2[20]) );
  DFFX1_RVT k2_reg_19_ ( .D(key[51]), .CLK(clk), .Q(k2[19]) );
  DFFX1_RVT k2_reg_18_ ( .D(key[50]), .CLK(clk), .Q(k2[18]) );
  DFFX1_RVT k2_reg_17_ ( .D(key[49]), .CLK(clk), .Q(k2[17]) );
  DFFX1_RVT k2_reg_16_ ( .D(key[48]), .CLK(clk), .Q(k2[16]) );
  DFFX1_RVT k2_reg_15_ ( .D(key[47]), .CLK(clk), .Q(k2[15]) );
  DFFX1_RVT k2_reg_14_ ( .D(key[46]), .CLK(clk), .Q(k2[14]) );
  DFFX1_RVT k2_reg_13_ ( .D(key[45]), .CLK(clk), .Q(k2[13]) );
  DFFX1_RVT k2_reg_12_ ( .D(key[44]), .CLK(clk), .Q(k2[12]) );
  DFFX1_RVT k2_reg_11_ ( .D(key[43]), .CLK(clk), .Q(k2[11]) );
  DFFX1_RVT k2_reg_10_ ( .D(key[42]), .CLK(clk), .Q(k2[10]) );
  DFFX1_RVT k2_reg_9_ ( .D(key[41]), .CLK(clk), .Q(k2[9]) );
  DFFX1_RVT k2_reg_8_ ( .D(key[40]), .CLK(clk), .Q(k2[8]) );
  DFFX1_RVT k2_reg_7_ ( .D(key[39]), .CLK(clk), .Q(k2[7]) );
  DFFX1_RVT k2_reg_6_ ( .D(key[38]), .CLK(clk), .Q(k2[6]) );
  DFFX1_RVT k2_reg_5_ ( .D(key[37]), .CLK(clk), .Q(k2[5]) );
  DFFX1_RVT k2_reg_4_ ( .D(key[36]), .CLK(clk), .Q(k2[4]) );
  DFFX1_RVT k2_reg_3_ ( .D(key[35]), .CLK(clk), .Q(k2[3]) );
  DFFX1_RVT k2_reg_2_ ( .D(key[34]), .CLK(clk), .Q(k2[2]) );
  DFFX1_RVT k2_reg_1_ ( .D(key[33]), .CLK(clk), .Q(k2[1]) );
  DFFX1_RVT k2_reg_0_ ( .D(key[32]), .CLK(clk), .Q(k2[0]) );
  DFFX1_RVT p03_reg_7_ ( .D(n1), .CLK(clk), .Q(p03[7]) );
  DFFX1_RVT p03_reg_6_ ( .D(n4), .CLK(clk), .Q(p03[6]) );
  DFFX1_RVT p03_reg_5_ ( .D(n5), .CLK(clk), .Q(p03[5]) );
  DFFX1_RVT p03_reg_4_ ( .D(n2), .CLK(clk), .Q(p03[4]) );
  DFFX1_RVT p03_reg_3_ ( .D(n7), .CLK(clk), .Q(p03[3]) );
  DFFX1_RVT p03_reg_2_ ( .D(n3), .CLK(clk), .Q(p03[2]) );
  DFFX1_RVT p03_reg_1_ ( .D(n6), .CLK(clk), .Q(p03[1]) );
  DFFX1_RVT p03_reg_0_ ( .D(n8), .CLK(clk), .Q(p03[0]) );
  INVX1_RVT U3 ( .A(n1842), .Y(n1) );
  INVX1_RVT U4 ( .A(n1594), .Y(n2) );
  INVX1_RVT U5 ( .A(n1405), .Y(n3) );
  INVX1_RVT U6 ( .A(n1765), .Y(n4) );
  INVX1_RVT U7 ( .A(n1674), .Y(n5) );
  INVX1_RVT U8 ( .A(n1180), .Y(n6) );
  INVX1_RVT U9 ( .A(n1503), .Y(n7) );
  INVX1_RVT U10 ( .A(n1066), .Y(n8) );
  INVX1_RVT U11 ( .A(n1580), .Y(n9) );
  INVX1_RVT U13 ( .A(n1569), .Y(n11) );
  INVX1_RVT U21 ( .A(n1697), .Y(n19) );
  INVX1_RVT U23 ( .A(n2582), .Y(n21) );
  INVX1_RVT U24 ( .A(n2334), .Y(n22) );
  INVX1_RVT U25 ( .A(n2145), .Y(n23) );
  INVX1_RVT U26 ( .A(n2505), .Y(n24) );
  INVX1_RVT U27 ( .A(n2414), .Y(n25) );
  INVX1_RVT U28 ( .A(n2039), .Y(n26) );
  INVX1_RVT U29 ( .A(n2243), .Y(n27) );
  INVX1_RVT U30 ( .A(n1925), .Y(n28) );
  INVX1_RVT U31 ( .A(n2320), .Y(n29) );
  INVX1_RVT U33 ( .A(n2309), .Y(n31) );
  INVX1_RVT U41 ( .A(n2437), .Y(n39) );
  INVX1_RVT U43 ( .A(n5022), .Y(n41) );
  INVX1_RVT U44 ( .A(n3074), .Y(n42) );
  INVX1_RVT U45 ( .A(n2885), .Y(n43) );
  INVX1_RVT U46 ( .A(n3902), .Y(n44) );
  INVX1_RVT U47 ( .A(n3154), .Y(n45) );
  INVX1_RVT U48 ( .A(n2779), .Y(n46) );
  INVX1_RVT U49 ( .A(n2983), .Y(n47) );
  INVX1_RVT U50 ( .A(n2665), .Y(n48) );
  INVX1_RVT U51 ( .A(n3060), .Y(n49) );
  INVX1_RVT U53 ( .A(n3049), .Y(n51) );
  INVX1_RVT U61 ( .A(n3177), .Y(n59) );
  INVX1_RVT U63 ( .A(n11996), .Y(n61) );
  INVX1_RVT U64 ( .A(n1286), .Y(n62) );
  INVX1_RVT U65 ( .A(n11007), .Y(n63) );
  INVX1_RVT U66 ( .A(n10017), .Y(n64) );
  INVX1_RVT U67 ( .A(n8044), .Y(n65) );
  INVX1_RVT U68 ( .A(n6954), .Y(n66) );
  INVX1_RVT U69 ( .A(n6114), .Y(n67) );
  INVX1_RVT U70 ( .A(n8875), .Y(n68) );
  INVX1_RVT U71 ( .A(n1361), .Y(n69) );
  INVX1_RVT U72 ( .A(n11056), .Y(n70) );
  INVX1_RVT U73 ( .A(n7034), .Y(n71) );
  INVX1_RVT U74 ( .A(n8901), .Y(n72) );
  INVX1_RVT U75 ( .A(n1312), .Y(n73) );
  INVX1_RVT U78 ( .A(n1328), .Y(n76) );
  INVX1_RVT U80 ( .A(n8065), .Y(n78) );
  INVX1_RVT U81 ( .A(n6131), .Y(n79) );
  INVX1_RVT U85 ( .A(n12014), .Y(n83) );
  INVX1_RVT U87 ( .A(n8063), .Y(n85) );
  INVX1_RVT U88 ( .A(n10435), .Y(n86) );
  INVX1_RVT U89 ( .A(n10187), .Y(n87) );
  INVX1_RVT U90 ( .A(n9919), .Y(n88) );
  INVX1_RVT U91 ( .A(n10358), .Y(n89) );
  INVX1_RVT U92 ( .A(n10267), .Y(n90) );
  INVX1_RVT U93 ( .A(n9813), .Y(n91) );
  INVX1_RVT U94 ( .A(n10096), .Y(n92) );
  INVX1_RVT U95 ( .A(n9699), .Y(n93) );
  INVX1_RVT U96 ( .A(n10173), .Y(n94) );
  INVX1_RVT U98 ( .A(n10162), .Y(n96) );
  INVX1_RVT U106 ( .A(n10290), .Y(n104) );
  INVX1_RVT U108 ( .A(n11256), .Y(n106) );
  INVX1_RVT U109 ( .A(n10927), .Y(n107) );
  INVX1_RVT U110 ( .A(n10738), .Y(n108) );
  INVX1_RVT U111 ( .A(n11179), .Y(n109) );
  INVX1_RVT U112 ( .A(n11088), .Y(n110) );
  INVX1_RVT U113 ( .A(n10632), .Y(n111) );
  INVX1_RVT U114 ( .A(n10836), .Y(n112) );
  INVX1_RVT U115 ( .A(n10518), .Y(n113) );
  INVX1_RVT U116 ( .A(n10913), .Y(n114) );
  INVX1_RVT U118 ( .A(n10902), .Y(n116) );
  INVX1_RVT U126 ( .A(n11111), .Y(n124) );
  INVX1_RVT U128 ( .A(n12066), .Y(n126) );
  INVX1_RVT U129 ( .A(n11748), .Y(n127) );
  INVX1_RVT U130 ( .A(n11559), .Y(n128) );
  INVX1_RVT U131 ( .A(n11919), .Y(n129) );
  INVX1_RVT U132 ( .A(n11828), .Y(n130) );
  INVX1_RVT U133 ( .A(n11453), .Y(n131) );
  INVX1_RVT U134 ( .A(n11657), .Y(n132) );
  INVX1_RVT U135 ( .A(n11339), .Y(n133) );
  INVX1_RVT U136 ( .A(n11734), .Y(n134) );
  INVX1_RVT U138 ( .A(n11723), .Y(n136) );
  INVX1_RVT U146 ( .A(n11851), .Y(n144) );
  INVX1_RVT U148 ( .A(n983), .Y(n146) );
  INVX1_RVT U149 ( .A(n735), .Y(n147) );
  INVX1_RVT U150 ( .A(n546), .Y(n148) );
  INVX1_RVT U151 ( .A(n906), .Y(n149) );
  INVX1_RVT U152 ( .A(n815), .Y(n150) );
  INVX1_RVT U153 ( .A(n440), .Y(n151) );
  INVX1_RVT U154 ( .A(n644), .Y(n152) );
  INVX1_RVT U155 ( .A(n326), .Y(n153) );
  INVX1_RVT U156 ( .A(n721), .Y(n154) );
  INVX1_RVT U158 ( .A(n710), .Y(n156) );
  INVX1_RVT U166 ( .A(n838), .Y(n164) );
  INVX1_RVT U168 ( .A(n7221), .Y(n166) );
  INVX1_RVT U169 ( .A(n6874), .Y(n167) );
  INVX1_RVT U170 ( .A(n6685), .Y(n168) );
  INVX1_RVT U171 ( .A(n7144), .Y(n169) );
  INVX1_RVT U172 ( .A(n7053), .Y(n170) );
  INVX1_RVT U173 ( .A(n6579), .Y(n171) );
  INVX1_RVT U174 ( .A(n6783), .Y(n172) );
  INVX1_RVT U175 ( .A(n6465), .Y(n173) );
  INVX1_RVT U176 ( .A(n6860), .Y(n174) );
  INVX1_RVT U178 ( .A(n6849), .Y(n176) );
  INVX1_RVT U186 ( .A(n7076), .Y(n184) );
  INVX1_RVT U188 ( .A(n7961), .Y(n186) );
  INVX1_RVT U189 ( .A(n7713), .Y(n187) );
  INVX1_RVT U190 ( .A(n7524), .Y(n188) );
  INVX1_RVT U191 ( .A(n7884), .Y(n189) );
  INVX1_RVT U192 ( .A(n7793), .Y(n190) );
  INVX1_RVT U193 ( .A(n7418), .Y(n191) );
  INVX1_RVT U194 ( .A(n7622), .Y(n192) );
  INVX1_RVT U195 ( .A(n7304), .Y(n193) );
  INVX1_RVT U196 ( .A(n7699), .Y(n194) );
  INVX1_RVT U198 ( .A(n7688), .Y(n196) );
  INVX1_RVT U206 ( .A(n7816), .Y(n204) );
  INVX1_RVT U208 ( .A(n8792), .Y(n206) );
  INVX1_RVT U209 ( .A(n8544), .Y(n207) );
  INVX1_RVT U210 ( .A(n8355), .Y(n208) );
  INVX1_RVT U211 ( .A(n8715), .Y(n209) );
  INVX1_RVT U212 ( .A(n8624), .Y(n210) );
  INVX1_RVT U213 ( .A(n8249), .Y(n211) );
  INVX1_RVT U214 ( .A(n8453), .Y(n212) );
  INVX1_RVT U215 ( .A(n8135), .Y(n213) );
  INVX1_RVT U216 ( .A(n8530), .Y(n214) );
  INVX1_RVT U218 ( .A(n8519), .Y(n216) );
  INVX1_RVT U226 ( .A(n8647), .Y(n224) );
  INVX1_RVT U228 ( .A(n9616), .Y(n226) );
  INVX1_RVT U229 ( .A(n9368), .Y(n227) );
  INVX1_RVT U230 ( .A(n9179), .Y(n228) );
  INVX1_RVT U231 ( .A(n9539), .Y(n229) );
  INVX1_RVT U232 ( .A(n9448), .Y(n230) );
  INVX1_RVT U233 ( .A(n9073), .Y(n231) );
  INVX1_RVT U234 ( .A(n9277), .Y(n232) );
  INVX1_RVT U235 ( .A(n8959), .Y(n233) );
  INVX1_RVT U236 ( .A(n9354), .Y(n234) );
  INVX1_RVT U238 ( .A(n9343), .Y(n236) );
  INVX1_RVT U246 ( .A(n9471), .Y(n244) );
  INVX1_RVT U248 ( .A(n3979), .Y(n246) );
  INVX1_RVT U249 ( .A(n3654), .Y(n247) );
  INVX1_RVT U250 ( .A(n3465), .Y(n248) );
  INVX1_RVT U251 ( .A(n3825), .Y(n249) );
  INVX1_RVT U252 ( .A(n3734), .Y(n250) );
  INVX1_RVT U253 ( .A(n3359), .Y(n251) );
  INVX1_RVT U254 ( .A(n3563), .Y(n252) );
  INVX1_RVT U255 ( .A(n3245), .Y(n253) );
  INVX1_RVT U256 ( .A(n3640), .Y(n254) );
  INVX1_RVT U258 ( .A(n3629), .Y(n256) );
  INVX1_RVT U266 ( .A(n3757), .Y(n264) );
  INVX1_RVT U268 ( .A(n4719), .Y(n266) );
  INVX1_RVT U269 ( .A(n4471), .Y(n267) );
  INVX1_RVT U270 ( .A(n4282), .Y(n268) );
  INVX1_RVT U271 ( .A(n4642), .Y(n269) );
  INVX1_RVT U272 ( .A(n4551), .Y(n270) );
  INVX1_RVT U273 ( .A(n4176), .Y(n271) );
  INVX1_RVT U274 ( .A(n4380), .Y(n272) );
  INVX1_RVT U275 ( .A(n4062), .Y(n273) );
  INVX1_RVT U276 ( .A(n4457), .Y(n274) );
  INVX1_RVT U278 ( .A(n4446), .Y(n276) );
  INVX1_RVT U286 ( .A(n4574), .Y(n284) );
  INVX1_RVT U288 ( .A(n5542), .Y(n286) );
  INVX1_RVT U289 ( .A(n5294), .Y(n287) );
  INVX1_RVT U290 ( .A(n5105), .Y(n288) );
  INVX1_RVT U291 ( .A(n5465), .Y(n289) );
  INVX1_RVT U292 ( .A(n5374), .Y(n290) );
  INVX1_RVT U293 ( .A(n4916), .Y(n291) );
  INVX1_RVT U294 ( .A(n5203), .Y(n292) );
  INVX1_RVT U295 ( .A(n4802), .Y(n293) );
  INVX1_RVT U296 ( .A(n5280), .Y(n294) );
  INVX1_RVT U298 ( .A(n5269), .Y(n296) );
  INVX1_RVT U306 ( .A(n5397), .Y(n304) );
  INVX1_RVT U308 ( .A(n6382), .Y(n306) );
  INVX1_RVT U309 ( .A(n6034), .Y(n307) );
  INVX1_RVT U310 ( .A(n5845), .Y(n308) );
  INVX1_RVT U311 ( .A(n6305), .Y(n309) );
  INVX1_RVT U312 ( .A(n6214), .Y(n310) );
  INVX1_RVT U313 ( .A(n5739), .Y(n311) );
  INVX1_RVT U314 ( .A(n5943), .Y(n312) );
  INVX1_RVT U315 ( .A(n5625), .Y(n313) );
  INVX1_RVT U316 ( .A(n6020), .Y(n314) );
  INVX1_RVT U318 ( .A(n6009), .Y(n316) );
  INVX1_RVT U326 ( .A(n6237), .Y(n324) );
  XOR2X1_RVT U328 ( .A1(p32[1]), .A2(k3[9]), .Y(out[9]) );
  XOR2X1_RVT U329 ( .A1(p03[3]), .A2(k0[3]), .Y(out[99]) );
  XOR2X1_RVT U330 ( .A1(p03[2]), .A2(k0[2]), .Y(out[98]) );
  XOR2X1_RVT U331 ( .A1(p03[1]), .A2(k0[1]), .Y(out[97]) );
  XOR2X1_RVT U332 ( .A1(p03[0]), .A2(k0[0]), .Y(out[96]) );
  XOR2X1_RVT U333 ( .A1(p10[7]), .A2(k1[31]), .Y(out[95]) );
  XOR2X1_RVT U334 ( .A1(p10[6]), .A2(k1[30]), .Y(out[94]) );
  XOR2X1_RVT U335 ( .A1(p10[5]), .A2(k1[29]), .Y(out[93]) );
  XOR2X1_RVT U336 ( .A1(p10[4]), .A2(k1[28]), .Y(out[92]) );
  XOR2X1_RVT U337 ( .A1(p10[3]), .A2(k1[27]), .Y(out[91]) );
  XOR2X1_RVT U338 ( .A1(p10[2]), .A2(k1[26]), .Y(out[90]) );
  XOR2X1_RVT U339 ( .A1(p32[0]), .A2(k3[8]), .Y(out[8]) );
  XOR2X1_RVT U340 ( .A1(p10[1]), .A2(k1[25]), .Y(out[89]) );
  XOR2X1_RVT U341 ( .A1(p10[0]), .A2(k1[24]), .Y(out[88]) );
  XOR2X1_RVT U342 ( .A1(p11[7]), .A2(k1[23]), .Y(out[87]) );
  XOR2X1_RVT U343 ( .A1(p11[6]), .A2(k1[22]), .Y(out[86]) );
  XOR2X1_RVT U344 ( .A1(p11[5]), .A2(k1[21]), .Y(out[85]) );
  XOR2X1_RVT U345 ( .A1(p11[4]), .A2(k1[20]), .Y(out[84]) );
  XOR2X1_RVT U346 ( .A1(p11[3]), .A2(k1[19]), .Y(out[83]) );
  XOR2X1_RVT U347 ( .A1(p11[2]), .A2(k1[18]), .Y(out[82]) );
  XOR2X1_RVT U348 ( .A1(p11[1]), .A2(k1[17]), .Y(out[81]) );
  XOR2X1_RVT U349 ( .A1(p11[0]), .A2(k1[16]), .Y(out[80]) );
  XOR2X1_RVT U350 ( .A1(p33[7]), .A2(k3[7]), .Y(out[7]) );
  XOR2X1_RVT U351 ( .A1(p12[7]), .A2(k1[15]), .Y(out[79]) );
  XOR2X1_RVT U352 ( .A1(p12[6]), .A2(k1[14]), .Y(out[78]) );
  XOR2X1_RVT U353 ( .A1(p12[5]), .A2(k1[13]), .Y(out[77]) );
  XOR2X1_RVT U354 ( .A1(p12[4]), .A2(k1[12]), .Y(out[76]) );
  XOR2X1_RVT U355 ( .A1(p12[3]), .A2(k1[11]), .Y(out[75]) );
  XOR2X1_RVT U356 ( .A1(p12[2]), .A2(k1[10]), .Y(out[74]) );
  XOR2X1_RVT U357 ( .A1(p12[1]), .A2(k1[9]), .Y(out[73]) );
  XOR2X1_RVT U358 ( .A1(p12[0]), .A2(k1[8]), .Y(out[72]) );
  XOR2X1_RVT U359 ( .A1(p13[7]), .A2(k1[7]), .Y(out[71]) );
  XOR2X1_RVT U360 ( .A1(p13[6]), .A2(k1[6]), .Y(out[70]) );
  XOR2X1_RVT U361 ( .A1(p33[6]), .A2(k3[6]), .Y(out[6]) );
  XOR2X1_RVT U362 ( .A1(p13[5]), .A2(k1[5]), .Y(out[69]) );
  XOR2X1_RVT U363 ( .A1(p13[4]), .A2(k1[4]), .Y(out[68]) );
  XOR2X1_RVT U364 ( .A1(p13[3]), .A2(k1[3]), .Y(out[67]) );
  XOR2X1_RVT U365 ( .A1(p13[2]), .A2(k1[2]), .Y(out[66]) );
  XOR2X1_RVT U366 ( .A1(p13[1]), .A2(k1[1]), .Y(out[65]) );
  XOR2X1_RVT U367 ( .A1(p13[0]), .A2(k1[0]), .Y(out[64]) );
  XOR2X1_RVT U368 ( .A1(p20[7]), .A2(k2[31]), .Y(out[63]) );
  XOR2X1_RVT U369 ( .A1(p20[6]), .A2(k2[30]), .Y(out[62]) );
  XOR2X1_RVT U370 ( .A1(p20[5]), .A2(k2[29]), .Y(out[61]) );
  XOR2X1_RVT U371 ( .A1(p20[4]), .A2(k2[28]), .Y(out[60]) );
  XOR2X1_RVT U372 ( .A1(p33[5]), .A2(k3[5]), .Y(out[5]) );
  XOR2X1_RVT U373 ( .A1(p20[3]), .A2(k2[27]), .Y(out[59]) );
  XOR2X1_RVT U374 ( .A1(p20[2]), .A2(k2[26]), .Y(out[58]) );
  XOR2X1_RVT U375 ( .A1(p20[1]), .A2(k2[25]), .Y(out[57]) );
  XOR2X1_RVT U376 ( .A1(p20[0]), .A2(k2[24]), .Y(out[56]) );
  XOR2X1_RVT U377 ( .A1(p21[7]), .A2(k2[23]), .Y(out[55]) );
  XOR2X1_RVT U378 ( .A1(p21[6]), .A2(k2[22]), .Y(out[54]) );
  XOR2X1_RVT U379 ( .A1(p21[5]), .A2(k2[21]), .Y(out[53]) );
  XOR2X1_RVT U380 ( .A1(p21[4]), .A2(k2[20]), .Y(out[52]) );
  XOR2X1_RVT U381 ( .A1(p21[3]), .A2(k2[19]), .Y(out[51]) );
  XOR2X1_RVT U382 ( .A1(p21[2]), .A2(k2[18]), .Y(out[50]) );
  XOR2X1_RVT U383 ( .A1(p33[4]), .A2(k3[4]), .Y(out[4]) );
  XOR2X1_RVT U384 ( .A1(p21[1]), .A2(k2[17]), .Y(out[49]) );
  XOR2X1_RVT U385 ( .A1(p21[0]), .A2(k2[16]), .Y(out[48]) );
  XOR2X1_RVT U386 ( .A1(p22[7]), .A2(k2[15]), .Y(out[47]) );
  XOR2X1_RVT U387 ( .A1(p22[6]), .A2(k2[14]), .Y(out[46]) );
  XOR2X1_RVT U388 ( .A1(p22[5]), .A2(k2[13]), .Y(out[45]) );
  XOR2X1_RVT U389 ( .A1(p22[4]), .A2(k2[12]), .Y(out[44]) );
  XOR2X1_RVT U390 ( .A1(p22[3]), .A2(k2[11]), .Y(out[43]) );
  XOR2X1_RVT U391 ( .A1(p22[2]), .A2(k2[10]), .Y(out[42]) );
  XOR2X1_RVT U392 ( .A1(p22[1]), .A2(k2[9]), .Y(out[41]) );
  XOR2X1_RVT U393 ( .A1(p22[0]), .A2(k2[8]), .Y(out[40]) );
  XOR2X1_RVT U394 ( .A1(p33[3]), .A2(k3[3]), .Y(out[3]) );
  XOR2X1_RVT U395 ( .A1(p23[7]), .A2(k2[7]), .Y(out[39]) );
  XOR2X1_RVT U396 ( .A1(p23[6]), .A2(k2[6]), .Y(out[38]) );
  XOR2X1_RVT U397 ( .A1(p23[5]), .A2(k2[5]), .Y(out[37]) );
  XOR2X1_RVT U398 ( .A1(p23[4]), .A2(k2[4]), .Y(out[36]) );
  XOR2X1_RVT U399 ( .A1(p23[3]), .A2(k2[3]), .Y(out[35]) );
  XOR2X1_RVT U400 ( .A1(p23[2]), .A2(k2[2]), .Y(out[34]) );
  XOR2X1_RVT U401 ( .A1(p23[1]), .A2(k2[1]), .Y(out[33]) );
  XOR2X1_RVT U402 ( .A1(p23[0]), .A2(k2[0]), .Y(out[32]) );
  XOR2X1_RVT U403 ( .A1(p30[7]), .A2(k3[31]), .Y(out[31]) );
  XOR2X1_RVT U404 ( .A1(p30[6]), .A2(k3[30]), .Y(out[30]) );
  XOR2X1_RVT U405 ( .A1(p33[2]), .A2(k3[2]), .Y(out[2]) );
  XOR2X1_RVT U406 ( .A1(p30[5]), .A2(k3[29]), .Y(out[29]) );
  XOR2X1_RVT U407 ( .A1(p30[4]), .A2(k3[28]), .Y(out[28]) );
  XOR2X1_RVT U408 ( .A1(p30[3]), .A2(k3[27]), .Y(out[27]) );
  XOR2X1_RVT U409 ( .A1(p30[2]), .A2(k3[26]), .Y(out[26]) );
  XOR2X1_RVT U410 ( .A1(p30[1]), .A2(k3[25]), .Y(out[25]) );
  XOR2X1_RVT U411 ( .A1(p30[0]), .A2(k3[24]), .Y(out[24]) );
  XOR2X1_RVT U412 ( .A1(p31[7]), .A2(k3[23]), .Y(out[23]) );
  XOR2X1_RVT U413 ( .A1(p31[6]), .A2(k3[22]), .Y(out[22]) );
  XOR2X1_RVT U414 ( .A1(p31[5]), .A2(k3[21]), .Y(out[21]) );
  XOR2X1_RVT U415 ( .A1(p31[4]), .A2(k3[20]), .Y(out[20]) );
  XOR2X1_RVT U416 ( .A1(p33[1]), .A2(k3[1]), .Y(out[1]) );
  XOR2X1_RVT U417 ( .A1(p31[3]), .A2(k3[19]), .Y(out[19]) );
  XOR2X1_RVT U418 ( .A1(p31[2]), .A2(k3[18]), .Y(out[18]) );
  XOR2X1_RVT U419 ( .A1(p31[1]), .A2(k3[17]), .Y(out[17]) );
  XOR2X1_RVT U420 ( .A1(p31[0]), .A2(k3[16]), .Y(out[16]) );
  XOR2X1_RVT U421 ( .A1(p32[7]), .A2(k3[15]), .Y(out[15]) );
  XOR2X1_RVT U422 ( .A1(p32[6]), .A2(k3[14]), .Y(out[14]) );
  XOR2X1_RVT U423 ( .A1(p32[5]), .A2(k3[13]), .Y(out[13]) );
  XOR2X1_RVT U424 ( .A1(p32[4]), .A2(k3[12]), .Y(out[12]) );
  XOR2X1_RVT U425 ( .A1(p00[7]), .A2(k0[31]), .Y(out[127]) );
  XOR2X1_RVT U426 ( .A1(p00[6]), .A2(k0[30]), .Y(out[126]) );
  XOR2X1_RVT U427 ( .A1(p00[5]), .A2(k0[29]), .Y(out[125]) );
  XOR2X1_RVT U428 ( .A1(p00[4]), .A2(k0[28]), .Y(out[124]) );
  XOR2X1_RVT U429 ( .A1(p00[3]), .A2(k0[27]), .Y(out[123]) );
  XOR2X1_RVT U430 ( .A1(p00[2]), .A2(k0[26]), .Y(out[122]) );
  XOR2X1_RVT U431 ( .A1(p00[1]), .A2(k0[25]), .Y(out[121]) );
  XOR2X1_RVT U432 ( .A1(p00[0]), .A2(k0[24]), .Y(out[120]) );
  XOR2X1_RVT U433 ( .A1(p32[3]), .A2(k3[11]), .Y(out[11]) );
  XOR2X1_RVT U434 ( .A1(p01[7]), .A2(k0[23]), .Y(out[119]) );
  XOR2X1_RVT U435 ( .A1(p01[6]), .A2(k0[22]), .Y(out[118]) );
  XOR2X1_RVT U436 ( .A1(p01[5]), .A2(k0[21]), .Y(out[117]) );
  XOR2X1_RVT U437 ( .A1(p01[4]), .A2(k0[20]), .Y(out[116]) );
  XOR2X1_RVT U438 ( .A1(p01[3]), .A2(k0[19]), .Y(out[115]) );
  XOR2X1_RVT U439 ( .A1(p01[2]), .A2(k0[18]), .Y(out[114]) );
  XOR2X1_RVT U440 ( .A1(p01[1]), .A2(k0[17]), .Y(out[113]) );
  XOR2X1_RVT U441 ( .A1(p01[0]), .A2(k0[16]), .Y(out[112]) );
  XOR2X1_RVT U442 ( .A1(p02[7]), .A2(k0[15]), .Y(out[111]) );
  XOR2X1_RVT U443 ( .A1(p02[6]), .A2(k0[14]), .Y(out[110]) );
  XOR2X1_RVT U444 ( .A1(p32[2]), .A2(k3[10]), .Y(out[10]) );
  XOR2X1_RVT U445 ( .A1(p02[5]), .A2(k0[13]), .Y(out[109]) );
  XOR2X1_RVT U446 ( .A1(p02[4]), .A2(k0[12]), .Y(out[108]) );
  XOR2X1_RVT U447 ( .A1(p02[3]), .A2(k0[11]), .Y(out[107]) );
  XOR2X1_RVT U448 ( .A1(p02[2]), .A2(k0[10]), .Y(out[106]) );
  XOR2X1_RVT U449 ( .A1(p02[1]), .A2(k0[9]), .Y(out[105]) );
  XOR2X1_RVT U450 ( .A1(p02[0]), .A2(k0[8]), .Y(out[104]) );
  XOR2X1_RVT U451 ( .A1(p03[7]), .A2(k0[7]), .Y(out[103]) );
  XOR2X1_RVT U452 ( .A1(p03[6]), .A2(k0[6]), .Y(out[102]) );
  XOR2X1_RVT U453 ( .A1(p03[5]), .A2(k0[5]), .Y(out[101]) );
  XOR2X1_RVT U454 ( .A1(p03[4]), .A2(k0[4]), .Y(out[100]) );
  XOR2X1_RVT U455 ( .A1(p33[0]), .A2(k3[0]), .Y(out[0]) );
  AND4X1_RVT U456 ( .A1(n327), .A2(n328), .A3(n329), .A4(n330), .Y(n326) );
  AND4X1_RVT U457 ( .A1(n331), .A2(n332), .A3(n333), .A4(n334), .Y(n330) );
  AND4X1_RVT U458 ( .A1(n335), .A2(n336), .A3(n337), .A4(n338), .Y(n334) );
  OR2X1_RVT U459 ( .A1(n12669), .A2(n340), .Y(n333) );
  OR2X1_RVT U460 ( .A1(n341), .A2(n342), .Y(n331) );
  OR2X1_RVT U461 ( .A1(n12816), .A2(n343), .Y(n342) );
  AND4X1_RVT U462 ( .A1(n344), .A2(n345), .A3(n346), .A4(n347), .Y(n329) );
  OR2X1_RVT U463 ( .A1(n348), .A2(n12814), .Y(n347) );
  AND2X1_RVT U464 ( .A1(n349), .A2(n350), .Y(n348) );
  AND2X1_RVT U465 ( .A1(n351), .A2(n352), .Y(n346) );
  OR2X1_RVT U466 ( .A1(n353), .A2(n156), .Y(n352) );
  AND2X1_RVT U467 ( .A1(n354), .A2(n355), .Y(n353) );
  OR2X1_RVT U468 ( .A1(n12660), .A2(n357), .Y(n355) );
  OR2X1_RVT U469 ( .A1(n343), .A2(n358), .Y(n354) );
  OR2X1_RVT U470 ( .A1(n359), .A2(n12666), .Y(n351) );
  AND2X1_RVT U471 ( .A1(n361), .A2(n362), .Y(n359) );
  OR2X1_RVT U472 ( .A1(n363), .A2(n364), .Y(n345) );
  AND2X1_RVT U473 ( .A1(n365), .A2(n366), .Y(n363) );
  OR2X1_RVT U474 ( .A1(n12661), .A2(n367), .Y(n366) );
  AND2X1_RVT U475 ( .A1(n368), .A2(n369), .Y(n365) );
  AND2X1_RVT U476 ( .A1(n370), .A2(n371), .Y(n344) );
  OR2X1_RVT U477 ( .A1(n372), .A2(n12643), .Y(n371) );
  AND2X1_RVT U478 ( .A1(n374), .A2(n375), .Y(n372) );
  OR2X1_RVT U479 ( .A1(n376), .A2(n377), .Y(n375) );
  OR2X1_RVT U480 ( .A1(n12652), .A2(n12647), .Y(n377) );
  OR2X1_RVT U481 ( .A1(n380), .A2(n381), .Y(n370) );
  AND2X1_RVT U482 ( .A1(n382), .A2(n383), .Y(n380) );
  AND2X1_RVT U483 ( .A1(n384), .A2(n385), .Y(n382) );
  AND4X1_RVT U484 ( .A1(n386), .A2(n387), .A3(n388), .A4(n389), .Y(n328) );
  AND4X1_RVT U485 ( .A1(n390), .A2(n391), .A3(n392), .A4(n393), .Y(n389) );
  OR2X1_RVT U486 ( .A1(n394), .A2(n12672), .Y(n393) );
  AND4X1_RVT U487 ( .A1(n396), .A2(n397), .A3(n398), .A4(n399), .Y(n394) );
  OR2X1_RVT U488 ( .A1(n400), .A2(n367), .Y(n399) );
  OR2X1_RVT U489 ( .A1(n401), .A2(n12658), .Y(n398) );
  OR2X1_RVT U490 ( .A1(n403), .A2(n12649), .Y(n392) );
  AND4X1_RVT U491 ( .A1(n404), .A2(n405), .A3(n406), .A4(n407), .Y(n403) );
  OR2X1_RVT U492 ( .A1(n408), .A2(n409), .Y(n407) );
  OR2X1_RVT U493 ( .A1(n12666), .A2(n12661), .Y(n409) );
  AND2X1_RVT U494 ( .A1(n410), .A2(n411), .Y(n406) );
  OR2X1_RVT U495 ( .A1(n12818), .A2(n412), .Y(n405) );
  OR2X1_RVT U496 ( .A1(n413), .A2(n414), .Y(n404) );
  AND2X1_RVT U497 ( .A1(n415), .A2(n416), .Y(n413) );
  OR2X1_RVT U498 ( .A1(n12666), .A2(n417), .Y(n416) );
  OR2X1_RVT U499 ( .A1(n350), .A2(n418), .Y(n391) );
  OR2X1_RVT U500 ( .A1(n417), .A2(n419), .Y(n390) );
  OR2X1_RVT U501 ( .A1(n420), .A2(n421), .Y(n388) );
  OR2X1_RVT U502 ( .A1(n422), .A2(n415), .Y(n387) );
  OR2X1_RVT U503 ( .A1(n423), .A2(n424), .Y(n386) );
  AND4X1_RVT U504 ( .A1(n425), .A2(n426), .A3(n427), .A4(n428), .Y(n327) );
  AND2X1_RVT U505 ( .A1(n429), .A2(n430), .Y(n428) );
  OR2X1_RVT U506 ( .A1(n414), .A2(n431), .Y(n430) );
  AND2X1_RVT U507 ( .A1(n432), .A2(n433), .Y(n429) );
  OR2X1_RVT U508 ( .A1(n434), .A2(n357), .Y(n433) );
  OR2X1_RVT U509 ( .A1(n358), .A2(n435), .Y(n432) );
  OR2X1_RVT U510 ( .A1(n154), .A2(n436), .Y(n427) );
  OR2X1_RVT U511 ( .A1(n437), .A2(n12656), .Y(n426) );
  OR2X1_RVT U512 ( .A1(n12659), .A2(n439), .Y(n425) );
  AND4X1_RVT U513 ( .A1(n441), .A2(n442), .A3(n443), .A4(n444), .Y(n440) );
  AND4X1_RVT U514 ( .A1(n445), .A2(n336), .A3(n446), .A4(n447), .Y(n444) );
  AND4X1_RVT U515 ( .A1(n448), .A2(n449), .A3(n450), .A4(n451), .Y(n447) );
  OR2X1_RVT U516 ( .A1(n357), .A2(n452), .Y(n451) );
  OR2X1_RVT U517 ( .A1(n453), .A2(n12671), .Y(n452) );
  OR2X1_RVT U518 ( .A1(n358), .A2(n454), .Y(n450) );
  OR2X1_RVT U519 ( .A1(n154), .A2(n12655), .Y(n454) );
  OR2X1_RVT U520 ( .A1(n455), .A2(n401), .Y(n449) );
  AND2X1_RVT U521 ( .A1(n412), .A2(n456), .Y(n455) );
  OR2X1_RVT U522 ( .A1(n457), .A2(n458), .Y(n448) );
  AND2X1_RVT U523 ( .A1(n459), .A2(n460), .Y(n457) );
  AND2X1_RVT U524 ( .A1(n461), .A2(n462), .Y(n446) );
  OR2X1_RVT U525 ( .A1(n408), .A2(n463), .Y(n462) );
  OR2X1_RVT U526 ( .A1(n464), .A2(n12816), .Y(n463) );
  OR2X1_RVT U527 ( .A1(n465), .A2(n466), .Y(n461) );
  OR2X1_RVT U528 ( .A1(n467), .A2(n12660), .Y(n466) );
  OR2X1_RVT U529 ( .A1(n343), .A2(n468), .Y(n336) );
  AND4X1_RVT U530 ( .A1(n469), .A2(n470), .A3(n471), .A4(n472), .Y(n443) );
  AND4X1_RVT U531 ( .A1(n473), .A2(n474), .A3(n475), .A4(n476), .Y(n472) );
  OR2X1_RVT U532 ( .A1(n477), .A2(n12674), .Y(n476) );
  AND2X1_RVT U533 ( .A1(n479), .A2(n480), .Y(n477) );
  OR2X1_RVT U534 ( .A1(n12643), .A2(n358), .Y(n480) );
  OR2X1_RVT U535 ( .A1(n481), .A2(n360), .Y(n475) );
  AND2X1_RVT U536 ( .A1(n482), .A2(n483), .Y(n481) );
  OR2X1_RVT U537 ( .A1(n484), .A2(n12815), .Y(n474) );
  AND2X1_RVT U538 ( .A1(n485), .A2(n486), .Y(n484) );
  OR2X1_RVT U539 ( .A1(n487), .A2(n436), .Y(n486) );
  AND2X1_RVT U540 ( .A1(n12674), .A2(n12658), .Y(n487) );
  OR2X1_RVT U541 ( .A1(n488), .A2(n12644), .Y(n473) );
  AND2X1_RVT U542 ( .A1(n490), .A2(n491), .Y(n488) );
  OR2X1_RVT U543 ( .A1(n492), .A2(n12650), .Y(n471) );
  AND2X1_RVT U544 ( .A1(n493), .A2(n494), .Y(n492) );
  OR2X1_RVT U545 ( .A1(n12658), .A2(n495), .Y(n494) );
  AND2X1_RVT U546 ( .A1(n496), .A2(n497), .Y(n493) );
  OR2X1_RVT U547 ( .A1(n498), .A2(n499), .Y(n496) );
  OR2X1_RVT U548 ( .A1(n343), .A2(n414), .Y(n499) );
  OR2X1_RVT U549 ( .A1(n500), .A2(n12812), .Y(n470) );
  AND2X1_RVT U550 ( .A1(n501), .A2(n502), .Y(n500) );
  OR2X1_RVT U551 ( .A1(n503), .A2(n504), .Y(n469) );
  AND2X1_RVT U552 ( .A1(n505), .A2(n506), .Y(n503) );
  AND2X1_RVT U553 ( .A1(n507), .A2(n508), .Y(n505) );
  OR2X1_RVT U554 ( .A1(n156), .A2(n436), .Y(n508) );
  OR2X1_RVT U555 ( .A1(n12668), .A2(n401), .Y(n507) );
  AND4X1_RVT U556 ( .A1(n509), .A2(n510), .A3(n511), .A4(n512), .Y(n442) );
  AND4X1_RVT U557 ( .A1(n513), .A2(n514), .A3(n515), .A4(n516), .Y(n512) );
  OR2X1_RVT U558 ( .A1(n436), .A2(n435), .Y(n516) );
  OR2X1_RVT U559 ( .A1(n367), .A2(n517), .Y(n515) );
  OR2X1_RVT U560 ( .A1(n400), .A2(n518), .Y(n514) );
  OR2X1_RVT U561 ( .A1(n343), .A2(n519), .Y(n513) );
  AND2X1_RVT U562 ( .A1(n520), .A2(n521), .Y(n511) );
  OR2X1_RVT U563 ( .A1(n12669), .A2(n522), .Y(n521) );
  OR2X1_RVT U564 ( .A1(n12648), .A2(n419), .Y(n520) );
  OR2X1_RVT U565 ( .A1(n523), .A2(n378), .Y(n510) );
  AND4X1_RVT U566 ( .A1(n524), .A2(n525), .A3(n526), .A4(n527), .Y(n523) );
  OR2X1_RVT U567 ( .A1(n528), .A2(n343), .Y(n526) );
  OR2X1_RVT U568 ( .A1(n12804), .A2(n529), .Y(n525) );
  OR2X1_RVT U569 ( .A1(n530), .A2(n12812), .Y(n524) );
  AND2X1_RVT U570 ( .A1(n421), .A2(n531), .Y(n530) );
  OR2X1_RVT U571 ( .A1(n423), .A2(n532), .Y(n509) );
  AND4X1_RVT U572 ( .A1(n533), .A2(n534), .A3(n535), .A4(n536), .Y(n441) );
  AND4X1_RVT U573 ( .A1(n537), .A2(n538), .A3(n539), .A4(n540), .Y(n536) );
  OR2X1_RVT U574 ( .A1(n12808), .A2(n541), .Y(n540) );
  OR2X1_RVT U575 ( .A1(n12809), .A2(n542), .Y(n539) );
  OR2X1_RVT U576 ( .A1(n12806), .A2(n543), .Y(n538) );
  OR2X1_RVT U577 ( .A1(n12642), .A2(n544), .Y(n537) );
  OR2X1_RVT U578 ( .A1(n545), .A2(n12649), .Y(n534) );
  AND4X1_RVT U579 ( .A1(n547), .A2(n548), .A3(n549), .A4(n550), .Y(n546) );
  AND4X1_RVT U580 ( .A1(n551), .A2(n552), .A3(n553), .A4(n554), .Y(n550) );
  AND4X1_RVT U581 ( .A1(n555), .A2(n332), .A3(n502), .A4(n556), .Y(n554) );
  OR2X1_RVT U582 ( .A1(n557), .A2(n12803), .Y(n332) );
  AND2X1_RVT U583 ( .A1(n558), .A2(n559), .Y(n557) );
  OR2X1_RVT U584 ( .A1(n376), .A2(n560), .Y(n559) );
  OR2X1_RVT U585 ( .A1(n561), .A2(n458), .Y(n558) );
  OR2X1_RVT U586 ( .A1(n562), .A2(n417), .Y(n555) );
  AND2X1_RVT U587 ( .A1(n563), .A2(n564), .Y(n562) );
  OR2X1_RVT U588 ( .A1(n12808), .A2(n401), .Y(n564) );
  OR2X1_RVT U589 ( .A1(n565), .A2(n360), .Y(n553) );
  AND2X1_RVT U590 ( .A1(n566), .A2(n567), .Y(n565) );
  OR2X1_RVT U591 ( .A1(n568), .A2(n12814), .Y(n567) );
  AND2X1_RVT U592 ( .A1(n408), .A2(n569), .Y(n568) );
  OR2X1_RVT U593 ( .A1(n570), .A2(n12669), .Y(n552) );
  AND2X1_RVT U594 ( .A1(n571), .A2(n572), .Y(n570) );
  OR2X1_RVT U595 ( .A1(n401), .A2(n367), .Y(n572) );
  OR2X1_RVT U596 ( .A1(n573), .A2(n12652), .Y(n551) );
  AND2X1_RVT U597 ( .A1(n485), .A2(n574), .Y(n573) );
  OR2X1_RVT U598 ( .A1(n414), .A2(n575), .Y(n485) );
  AND4X1_RVT U599 ( .A1(n576), .A2(n577), .A3(n578), .A4(n579), .Y(n549) );
  OR2X1_RVT U600 ( .A1(n580), .A2(n12659), .Y(n579) );
  AND2X1_RVT U601 ( .A1(n581), .A2(n582), .Y(n580) );
  OR2X1_RVT U602 ( .A1(n458), .A2(n358), .Y(n582) );
  AND2X1_RVT U603 ( .A1(n583), .A2(n584), .Y(n581) );
  OR2X1_RVT U604 ( .A1(n498), .A2(n560), .Y(n583) );
  AND2X1_RVT U605 ( .A1(n585), .A2(n586), .Y(n578) );
  OR2X1_RVT U606 ( .A1(n587), .A2(n489), .Y(n586) );
  AND2X1_RVT U607 ( .A1(n588), .A2(n397), .Y(n587) );
  OR2X1_RVT U608 ( .A1(n343), .A2(n458), .Y(n397) );
  OR2X1_RVT U609 ( .A1(n589), .A2(n156), .Y(n585) );
  AND2X1_RVT U610 ( .A1(n590), .A2(n591), .Y(n589) );
  OR2X1_RVT U611 ( .A1(n592), .A2(n12661), .Y(n591) );
  AND2X1_RVT U612 ( .A1(n593), .A2(n594), .Y(n592) );
  OR2X1_RVT U613 ( .A1(n12656), .A2(n408), .Y(n594) );
  OR2X1_RVT U614 ( .A1(n12818), .A2(n12658), .Y(n593) );
  AND2X1_RVT U615 ( .A1(n459), .A2(n569), .Y(n590) );
  OR2X1_RVT U616 ( .A1(n489), .A2(n595), .Y(n459) );
  OR2X1_RVT U617 ( .A1(n12813), .A2(n12809), .Y(n595) );
  OR2X1_RVT U618 ( .A1(n596), .A2(n478), .Y(n577) );
  AND4X1_RVT U619 ( .A1(n437), .A2(n597), .A3(n598), .A4(n599), .Y(n596) );
  OR2X1_RVT U620 ( .A1(n12660), .A2(n458), .Y(n599) );
  AND2X1_RVT U621 ( .A1(n600), .A2(n601), .Y(n598) );
  OR2X1_RVT U622 ( .A1(n12818), .A2(n12669), .Y(n597) );
  AND2X1_RVT U623 ( .A1(n602), .A2(n603), .Y(n437) );
  OR2X1_RVT U624 ( .A1(n604), .A2(n154), .Y(n603) );
  OR2X1_RVT U625 ( .A1(n401), .A2(n12803), .Y(n602) );
  AND2X1_RVT U626 ( .A1(n605), .A2(n606), .Y(n576) );
  OR2X1_RVT U627 ( .A1(n607), .A2(n12805), .Y(n606) );
  AND2X1_RVT U628 ( .A1(n608), .A2(n609), .Y(n607) );
  OR2X1_RVT U629 ( .A1(n610), .A2(n12663), .Y(n609) );
  AND2X1_RVT U630 ( .A1(n611), .A2(n612), .Y(n610) );
  AND2X1_RVT U631 ( .A1(n613), .A2(n614), .Y(n608) );
  OR2X1_RVT U632 ( .A1(n615), .A2(n12672), .Y(n605) );
  AND4X1_RVT U633 ( .A1(n616), .A2(n617), .A3(n618), .A4(n619), .Y(n615) );
  OR2X1_RVT U634 ( .A1(n12817), .A2(n620), .Y(n618) );
  OR2X1_RVT U635 ( .A1(n154), .A2(n415), .Y(n617) );
  OR2X1_RVT U636 ( .A1(n504), .A2(n458), .Y(n616) );
  AND4X1_RVT U637 ( .A1(n621), .A2(n622), .A3(n623), .A4(n624), .Y(n548) );
  AND2X1_RVT U638 ( .A1(n625), .A2(n468), .Y(n624) );
  OR2X1_RVT U639 ( .A1(n12647), .A2(n434), .Y(n468) );
  AND2X1_RVT U640 ( .A1(n626), .A2(n627), .Y(n625) );
  OR2X1_RVT U641 ( .A1(n628), .A2(n383), .Y(n627) );
  OR2X1_RVT U642 ( .A1(n435), .A2(n495), .Y(n626) );
  OR2X1_RVT U643 ( .A1(n154), .A2(n629), .Y(n623) );
  OR2X1_RVT U644 ( .A1(n12816), .A2(n630), .Y(n622) );
  OR2X1_RVT U645 ( .A1(n504), .A2(n631), .Y(n621) );
  AND4X1_RVT U646 ( .A1(n632), .A2(n633), .A3(n634), .A4(n635), .Y(n547) );
  AND2X1_RVT U647 ( .A1(n636), .A2(n637), .Y(n635) );
  OR2X1_RVT U648 ( .A1(n12642), .A2(n638), .Y(n637) );
  AND2X1_RVT U649 ( .A1(n639), .A2(n640), .Y(n636) );
  OR2X1_RVT U650 ( .A1(n400), .A2(n410), .Y(n640) );
  OR2X1_RVT U651 ( .A1(n12663), .A2(n460), .Y(n410) );
  OR2X1_RVT U652 ( .A1(n12649), .A2(n641), .Y(n639) );
  OR2X1_RVT U653 ( .A1(n381), .A2(n374), .Y(n634) );
  OR2X1_RVT U654 ( .A1(n467), .A2(n642), .Y(n374) );
  OR2X1_RVT U655 ( .A1(n12812), .A2(n643), .Y(n633) );
  OR2X1_RVT U656 ( .A1(n12661), .A2(n501), .Y(n632) );
  OR2X1_RVT U657 ( .A1(n12803), .A2(n563), .Y(n501) );
  AND4X1_RVT U658 ( .A1(n645), .A2(n646), .A3(n647), .A4(n648), .Y(n644) );
  AND4X1_RVT U659 ( .A1(n649), .A2(n650), .A3(n651), .A4(n652), .Y(n648) );
  OR2X1_RVT U660 ( .A1(n164), .A2(n653), .Y(n652) );
  OR2X1_RVT U661 ( .A1(n654), .A2(n12674), .Y(n653) );
  AND2X1_RVT U662 ( .A1(n12663), .A2(n420), .Y(n654) );
  AND2X1_RVT U663 ( .A1(n335), .A2(n655), .Y(n651) );
  OR2X1_RVT U664 ( .A1(n12652), .A2(n656), .Y(n335) );
  OR2X1_RVT U665 ( .A1(n164), .A2(n414), .Y(n656) );
  OR2X1_RVT U666 ( .A1(n657), .A2(n343), .Y(n650) );
  AND2X1_RVT U667 ( .A1(n658), .A2(n659), .Y(n657) );
  AND2X1_RVT U668 ( .A1(n660), .A2(n661), .Y(n649) );
  OR2X1_RVT U669 ( .A1(n662), .A2(n663), .Y(n661) );
  AND2X1_RVT U670 ( .A1(n664), .A2(n424), .Y(n662) );
  OR2X1_RVT U671 ( .A1(n665), .A2(n415), .Y(n660) );
  AND2X1_RVT U672 ( .A1(n600), .A2(n434), .Y(n665) );
  OR2X1_RVT U673 ( .A1(n12650), .A2(n666), .Y(n600) );
  OR2X1_RVT U674 ( .A1(n12818), .A2(n12660), .Y(n666) );
  AND4X1_RVT U675 ( .A1(n667), .A2(n668), .A3(n669), .A4(n670), .Y(n647) );
  OR2X1_RVT U676 ( .A1(n671), .A2(n12808), .Y(n670) );
  AND2X1_RVT U677 ( .A1(n483), .A2(n672), .Y(n671) );
  OR2X1_RVT U678 ( .A1(n12816), .A2(n528), .Y(n483) );
  AND2X1_RVT U679 ( .A1(n673), .A2(n674), .Y(n669) );
  OR2X1_RVT U680 ( .A1(n675), .A2(n12806), .Y(n674) );
  AND2X1_RVT U681 ( .A1(n676), .A2(n677), .Y(n675) );
  OR2X1_RVT U682 ( .A1(n378), .A2(n620), .Y(n677) );
  OR2X1_RVT U683 ( .A1(n678), .A2(n12804), .Y(n673) );
  AND2X1_RVT U684 ( .A1(n679), .A2(n680), .Y(n678) );
  OR2X1_RVT U685 ( .A1(n681), .A2(n12663), .Y(n668) );
  AND2X1_RVT U686 ( .A1(n682), .A2(n683), .Y(n681) );
  AND2X1_RVT U687 ( .A1(n684), .A2(n685), .Y(n682) );
  AND2X1_RVT U688 ( .A1(n686), .A2(n687), .Y(n667) );
  OR2X1_RVT U689 ( .A1(n688), .A2(n604), .Y(n687) );
  AND2X1_RVT U690 ( .A1(n689), .A2(n435), .Y(n688) );
  AND2X1_RVT U691 ( .A1(n690), .A2(n691), .Y(n689) );
  OR2X1_RVT U692 ( .A1(n692), .A2(n12666), .Y(n686) );
  AND2X1_RVT U693 ( .A1(n693), .A2(n694), .Y(n692) );
  OR2X1_RVT U694 ( .A1(n12815), .A2(n12668), .Y(n694) );
  AND2X1_RVT U695 ( .A1(n424), .A2(n695), .Y(n693) );
  AND4X1_RVT U696 ( .A1(n696), .A2(n697), .A3(n698), .A4(n699), .Y(n646) );
  AND2X1_RVT U697 ( .A1(n700), .A2(n701), .Y(n699) );
  OR2X1_RVT U698 ( .A1(n417), .A2(n491), .Y(n701) );
  OR2X1_RVT U699 ( .A1(n12810), .A2(n424), .Y(n491) );
  AND2X1_RVT U700 ( .A1(n702), .A2(n703), .Y(n700) );
  OR2X1_RVT U701 ( .A1(n569), .A2(n383), .Y(n703) );
  OR2X1_RVT U702 ( .A1(n12817), .A2(n12659), .Y(n383) );
  OR2X1_RVT U703 ( .A1(n467), .A2(n517), .Y(n702) );
  OR2X1_RVT U704 ( .A1(n12805), .A2(n704), .Y(n517) );
  OR2X1_RVT U705 ( .A1(n705), .A2(n12642), .Y(n698) );
  AND4X1_RVT U706 ( .A1(n706), .A2(n707), .A3(n708), .A4(n709), .Y(n705) );
  OR2X1_RVT U707 ( .A1(n642), .A2(n415), .Y(n708) );
  OR2X1_RVT U708 ( .A1(n710), .A2(n412), .Y(n707) );
  OR2X1_RVT U709 ( .A1(n12814), .A2(n367), .Y(n706) );
  OR2X1_RVT U710 ( .A1(n711), .A2(n12643), .Y(n697) );
  AND2X1_RVT U711 ( .A1(n712), .A2(n713), .Y(n711) );
  OR2X1_RVT U712 ( .A1(n642), .A2(n367), .Y(n713) );
  AND2X1_RVT U713 ( .A1(n714), .A2(n643), .Y(n712) );
  OR2X1_RVT U714 ( .A1(n415), .A2(n715), .Y(n643) );
  OR2X1_RVT U715 ( .A1(n12805), .A2(n12817), .Y(n715) );
  OR2X1_RVT U716 ( .A1(n716), .A2(n12650), .Y(n696) );
  AND4X1_RVT U717 ( .A1(n717), .A2(n630), .A3(n439), .A4(n411), .Y(n716) );
  OR2X1_RVT U718 ( .A1(n436), .A2(n718), .Y(n411) );
  OR2X1_RVT U719 ( .A1(n12807), .A2(n373), .Y(n718) );
  OR2X1_RVT U720 ( .A1(n498), .A2(n532), .Y(n439) );
  OR2X1_RVT U721 ( .A1(n417), .A2(n719), .Y(n630) );
  OR2X1_RVT U722 ( .A1(n12674), .A2(n12643), .Y(n719) );
  OR2X1_RVT U723 ( .A1(n376), .A2(n720), .Y(n717) );
  OR2X1_RVT U724 ( .A1(n721), .A2(n12648), .Y(n720) );
  AND4X1_RVT U725 ( .A1(n722), .A2(n723), .A3(n724), .A4(n725), .Y(n645) );
  AND2X1_RVT U726 ( .A1(n726), .A2(n727), .Y(n725) );
  AND2X1_RVT U727 ( .A1(n728), .A2(n729), .Y(n726) );
  OR2X1_RVT U728 ( .A1(n408), .A2(n683), .Y(n729) );
  OR2X1_RVT U729 ( .A1(n420), .A2(n730), .Y(n683) );
  OR2X1_RVT U730 ( .A1(n12806), .A2(n12808), .Y(n730) );
  OR2X1_RVT U731 ( .A1(n12813), .A2(n731), .Y(n728) );
  OR2X1_RVT U732 ( .A1(n12659), .A2(n732), .Y(n724) );
  OR2X1_RVT U733 ( .A1(n12816), .A2(n733), .Y(n723) );
  OR2X1_RVT U734 ( .A1(n420), .A2(n734), .Y(n722) );
  AND4X1_RVT U735 ( .A1(n736), .A2(n737), .A3(n738), .A4(n739), .Y(n735) );
  AND4X1_RVT U736 ( .A1(n740), .A2(n741), .A3(n742), .A4(n743), .Y(n739) );
  AND4X1_RVT U737 ( .A1(n744), .A2(n745), .A3(n337), .A4(n746), .Y(n743) );
  OR2X1_RVT U738 ( .A1(n478), .A2(n747), .Y(n337) );
  OR2X1_RVT U739 ( .A1(n569), .A2(n156), .Y(n747) );
  OR2X1_RVT U740 ( .A1(n341), .A2(n748), .Y(n745) );
  OR2X1_RVT U741 ( .A1(n12811), .A2(n12814), .Y(n748) );
  OR2X1_RVT U742 ( .A1(n604), .A2(n749), .Y(n744) );
  OR2X1_RVT U743 ( .A1(n750), .A2(n378), .Y(n749) );
  AND2X1_RVT U744 ( .A1(n12663), .A2(n478), .Y(n750) );
  OR2X1_RVT U745 ( .A1(n751), .A2(n12669), .Y(n742) );
  AND2X1_RVT U746 ( .A1(n619), .A2(n691), .Y(n751) );
  OR2X1_RVT U747 ( .A1(n156), .A2(n752), .Y(n691) );
  OR2X1_RVT U748 ( .A1(n12642), .A2(n12810), .Y(n752) );
  OR2X1_RVT U749 ( .A1(n408), .A2(n753), .Y(n619) );
  OR2X1_RVT U750 ( .A1(n12808), .A2(n400), .Y(n753) );
  OR2X1_RVT U751 ( .A1(n754), .A2(n358), .Y(n741) );
  AND2X1_RVT U752 ( .A1(n755), .A2(n563), .Y(n754) );
  OR2X1_RVT U753 ( .A1(n464), .A2(n458), .Y(n740) );
  AND4X1_RVT U754 ( .A1(n756), .A2(n757), .A3(n758), .A4(n759), .Y(n738) );
  AND2X1_RVT U755 ( .A1(n760), .A2(n761), .Y(n759) );
  OR2X1_RVT U756 ( .A1(n762), .A2(n12663), .Y(n761) );
  AND2X1_RVT U757 ( .A1(n763), .A2(n431), .Y(n762) );
  AND2X1_RVT U758 ( .A1(n764), .A2(n765), .Y(n760) );
  OR2X1_RVT U759 ( .A1(n766), .A2(n414), .Y(n765) );
  AND2X1_RVT U760 ( .A1(n385), .A2(n357), .Y(n766) );
  OR2X1_RVT U761 ( .A1(n12816), .A2(n456), .Y(n385) );
  OR2X1_RVT U762 ( .A1(n767), .A2(n467), .Y(n764) );
  AND2X1_RVT U763 ( .A1(n659), .A2(n768), .Y(n767) );
  OR2X1_RVT U764 ( .A1(n12817), .A2(n495), .Y(n659) );
  OR2X1_RVT U765 ( .A1(n769), .A2(n12808), .Y(n758) );
  AND2X1_RVT U766 ( .A1(n362), .A2(n770), .Y(n769) );
  OR2X1_RVT U767 ( .A1(n498), .A2(n422), .Y(n770) );
  OR2X1_RVT U768 ( .A1(n401), .A2(n604), .Y(n362) );
  OR2X1_RVT U769 ( .A1(n771), .A2(n154), .Y(n757) );
  AND2X1_RVT U770 ( .A1(n412), .A2(n772), .Y(n771) );
  OR2X1_RVT U771 ( .A1(n773), .A2(n12647), .Y(n772) );
  AND2X1_RVT U772 ( .A1(n774), .A2(n775), .Y(n773) );
  OR2X1_RVT U773 ( .A1(n12809), .A2(n395), .Y(n775) );
  OR2X1_RVT U774 ( .A1(n12674), .A2(n498), .Y(n412) );
  OR2X1_RVT U775 ( .A1(n776), .A2(n482), .Y(n756) );
  AND2X1_RVT U776 ( .A1(n415), .A2(n460), .Y(n776) );
  OR2X1_RVT U777 ( .A1(n12805), .A2(n343), .Y(n460) );
  AND4X1_RVT U778 ( .A1(n777), .A2(n778), .A3(n779), .A4(n780), .Y(n737) );
  AND4X1_RVT U779 ( .A1(n781), .A2(n782), .A3(n783), .A4(n784), .Y(n780) );
  OR2X1_RVT U780 ( .A1(n785), .A2(n12816), .Y(n784) );
  AND2X1_RVT U781 ( .A1(n518), .A2(n786), .Y(n785) );
  OR2X1_RVT U782 ( .A1(n12671), .A2(n367), .Y(n786) );
  OR2X1_RVT U783 ( .A1(n787), .A2(n360), .Y(n783) );
  AND2X1_RVT U784 ( .A1(n788), .A2(n789), .Y(n787) );
  OR2X1_RVT U785 ( .A1(n790), .A2(n395), .Y(n789) );
  AND2X1_RVT U786 ( .A1(n420), .A2(n408), .Y(n790) );
  AND2X1_RVT U787 ( .A1(n422), .A2(n664), .Y(n788) );
  OR2X1_RVT U788 ( .A1(n12672), .A2(n560), .Y(n664) );
  OR2X1_RVT U789 ( .A1(n791), .A2(n12661), .Y(n782) );
  AND2X1_RVT U790 ( .A1(n792), .A2(n793), .Y(n791) );
  OR2X1_RVT U791 ( .A1(n408), .A2(n794), .Y(n793) );
  AND2X1_RVT U792 ( .A1(n490), .A2(n684), .Y(n792) );
  OR2X1_RVT U793 ( .A1(n400), .A2(n575), .Y(n684) );
  OR2X1_RVT U794 ( .A1(n373), .A2(n795), .Y(n490) );
  OR2X1_RVT U795 ( .A1(n796), .A2(n343), .Y(n781) );
  AND4X1_RVT U796 ( .A1(n797), .A2(n798), .A3(n799), .A4(n732), .Y(n796) );
  OR2X1_RVT U797 ( .A1(n436), .A2(n800), .Y(n732) );
  OR2X1_RVT U798 ( .A1(n12642), .A2(n400), .Y(n800) );
  OR2X1_RVT U799 ( .A1(n12813), .A2(n642), .Y(n798) );
  OR2X1_RVT U800 ( .A1(n401), .A2(n498), .Y(n797) );
  OR2X1_RVT U801 ( .A1(n569), .A2(n611), .Y(n779) );
  OR2X1_RVT U802 ( .A1(n801), .A2(n12645), .Y(n778) );
  AND4X1_RVT U803 ( .A1(n802), .A2(n803), .A3(n445), .A4(n543), .Y(n801) );
  OR2X1_RVT U804 ( .A1(n367), .A2(n532), .Y(n543) );
  OR2X1_RVT U805 ( .A1(n12813), .A2(n154), .Y(n532) );
  OR2X1_RVT U806 ( .A1(n360), .A2(n424), .Y(n445) );
  OR2X1_RVT U807 ( .A1(n12805), .A2(n795), .Y(n777) );
  AND4X1_RVT U808 ( .A1(n804), .A2(n805), .A3(n806), .A4(n807), .Y(n736) );
  OR2X1_RVT U809 ( .A1(n12650), .A2(n808), .Y(n807) );
  AND2X1_RVT U810 ( .A1(n809), .A2(n810), .Y(n806) );
  OR2X1_RVT U811 ( .A1(n12671), .A2(n563), .Y(n810) );
  OR2X1_RVT U812 ( .A1(n350), .A2(n424), .Y(n809) );
  OR2X1_RVT U813 ( .A1(n156), .A2(n381), .Y(n424) );
  OR2X1_RVT U814 ( .A1(n12674), .A2(n542), .Y(n805) );
  OR2X1_RVT U815 ( .A1(n417), .A2(n811), .Y(n542) );
  AND2X1_RVT U816 ( .A1(n812), .A2(n813), .Y(n804) );
  OR2X1_RVT U817 ( .A1(n12643), .A2(n814), .Y(n813) );
  OR2X1_RVT U818 ( .A1(n420), .A2(n369), .Y(n812) );
  OR2X1_RVT U819 ( .A1(n343), .A2(n628), .Y(n369) );
  AND4X1_RVT U820 ( .A1(n816), .A2(n817), .A3(n818), .A4(n819), .Y(n815) );
  AND4X1_RVT U821 ( .A1(n820), .A2(n821), .A3(n822), .A4(n823), .Y(n819) );
  AND4X1_RVT U822 ( .A1(n556), .A2(n746), .A3(n824), .A4(n825), .Y(n823) );
  OR2X1_RVT U823 ( .A1(n826), .A2(n827), .Y(n746) );
  OR2X1_RVT U824 ( .A1(n341), .A2(n611), .Y(n556) );
  OR2X1_RVT U825 ( .A1(n12814), .A2(n12659), .Y(n611) );
  AND4X1_RVT U826 ( .A1(n814), .A2(n680), .A3(n803), .A4(n338), .Y(n822) );
  OR2X1_RVT U827 ( .A1(n828), .A2(n528), .Y(n338) );
  OR2X1_RVT U828 ( .A1(n343), .A2(n829), .Y(n803) );
  OR2X1_RVT U829 ( .A1(n376), .A2(n154), .Y(n680) );
  OR2X1_RVT U830 ( .A1(n367), .A2(n830), .Y(n814) );
  OR2X1_RVT U831 ( .A1(n12649), .A2(n12669), .Y(n830) );
  AND4X1_RVT U832 ( .A1(n831), .A2(n832), .A3(n833), .A4(n834), .Y(n821) );
  OR2X1_RVT U833 ( .A1(n620), .A2(n835), .Y(n834) );
  OR2X1_RVT U834 ( .A1(n12669), .A2(n400), .Y(n835) );
  OR2X1_RVT U835 ( .A1(n529), .A2(n836), .Y(n833) );
  OR2X1_RVT U836 ( .A1(n12815), .A2(n417), .Y(n836) );
  OR2X1_RVT U837 ( .A1(n755), .A2(n837), .Y(n832) );
  OR2X1_RVT U838 ( .A1(n838), .A2(n414), .Y(n837) );
  OR2X1_RVT U839 ( .A1(n12666), .A2(n839), .Y(n831) );
  OR2X1_RVT U840 ( .A1(n840), .A2(n12649), .Y(n839) );
  AND2X1_RVT U841 ( .A1(n628), .A2(n841), .Y(n840) );
  AND2X1_RVT U842 ( .A1(n842), .A2(n843), .Y(n820) );
  OR2X1_RVT U843 ( .A1(n844), .A2(n395), .Y(n843) );
  AND2X1_RVT U844 ( .A1(n845), .A2(n846), .Y(n844) );
  OR2X1_RVT U845 ( .A1(n12648), .A2(n588), .Y(n846) );
  OR2X1_RVT U846 ( .A1(n12652), .A2(n663), .Y(n845) );
  AND2X1_RVT U847 ( .A1(n847), .A2(n848), .Y(n842) );
  OR2X1_RVT U848 ( .A1(n849), .A2(n434), .Y(n848) );
  AND2X1_RVT U849 ( .A1(n850), .A2(n851), .Y(n849) );
  OR2X1_RVT U850 ( .A1(n12655), .A2(n164), .Y(n851) );
  NAND2X1_RVT U851 ( .A1(n417), .A2(n12807), .Y(n850) );
  OR2X1_RVT U852 ( .A1(n852), .A2(n156), .Y(n847) );
  AND2X1_RVT U853 ( .A1(n641), .A2(n518), .Y(n852) );
  OR2X1_RVT U854 ( .A1(n367), .A2(n853), .Y(n518) );
  OR2X1_RVT U855 ( .A1(n12818), .A2(n12644), .Y(n853) );
  AND4X1_RVT U856 ( .A1(n535), .A2(n854), .A3(n727), .A4(n855), .Y(n818) );
  AND4X1_RVT U857 ( .A1(n856), .A2(n857), .A3(n858), .A4(n859), .Y(n855) );
  OR2X1_RVT U858 ( .A1(n498), .A2(n419), .Y(n859) );
  OR2X1_RVT U859 ( .A1(n436), .A2(n465), .Y(n858) );
  OR2X1_RVT U860 ( .A1(n12806), .A2(n690), .Y(n857) );
  OR2X1_RVT U861 ( .A1(n414), .A2(n396), .Y(n690) );
  OR2X1_RVT U862 ( .A1(n12814), .A2(n478), .Y(n396) );
  OR2X1_RVT U863 ( .A1(n12658), .A2(n519), .Y(n856) );
  OR2X1_RVT U864 ( .A1(n400), .A2(n628), .Y(n519) );
  OR2X1_RVT U865 ( .A1(n12642), .A2(n604), .Y(n628) );
  AND2X1_RVT U866 ( .A1(n860), .A2(n861), .Y(n727) );
  OR2X1_RVT U867 ( .A1(n862), .A2(n467), .Y(n861) );
  OR2X1_RVT U868 ( .A1(n12668), .A2(n156), .Y(n862) );
  OR2X1_RVT U869 ( .A1(n863), .A2(n350), .Y(n860) );
  OR2X1_RVT U870 ( .A1(n12805), .A2(n467), .Y(n350) );
  OR2X1_RVT U871 ( .A1(n364), .A2(n414), .Y(n863) );
  OR2X1_RVT U872 ( .A1(n12650), .A2(n733), .Y(n854) );
  AND2X1_RVT U873 ( .A1(n864), .A2(n865), .Y(n535) );
  OR2X1_RVT U874 ( .A1(n418), .A2(n456), .Y(n865) );
  OR2X1_RVT U875 ( .A1(n866), .A2(n867), .Y(n864) );
  AND4X1_RVT U876 ( .A1(n868), .A2(n869), .A3(n870), .A4(n871), .Y(n817) );
  OR2X1_RVT U877 ( .A1(n872), .A2(n604), .Y(n871) );
  AND2X1_RVT U878 ( .A1(n873), .A2(n613), .Y(n872) );
  OR2X1_RVT U879 ( .A1(n12656), .A2(n829), .Y(n613) );
  OR2X1_RVT U880 ( .A1(n874), .A2(n12811), .Y(n870) );
  AND2X1_RVT U881 ( .A1(n541), .A2(n506), .Y(n874) );
  OR2X1_RVT U882 ( .A1(n12805), .A2(n482), .Y(n506) );
  OR2X1_RVT U883 ( .A1(n875), .A2(n561), .Y(n869) );
  AND2X1_RVT U884 ( .A1(n876), .A2(n877), .Y(n875) );
  OR2X1_RVT U885 ( .A1(n12645), .A2(n420), .Y(n877) );
  AND2X1_RVT U886 ( .A1(n878), .A2(n458), .Y(n876) );
  OR2X1_RVT U887 ( .A1(n154), .A2(n417), .Y(n878) );
  OR2X1_RVT U888 ( .A1(n879), .A2(n358), .Y(n868) );
  AND2X1_RVT U889 ( .A1(n880), .A2(n881), .Y(n879) );
  NAND2X1_RVT U890 ( .A1(n343), .A2(n721), .Y(n881) );
  AND2X1_RVT U891 ( .A1(n882), .A2(n571), .Y(n880) );
  OR2X1_RVT U892 ( .A1(n504), .A2(n829), .Y(n571) );
  OR2X1_RVT U893 ( .A1(n12665), .A2(n883), .Y(n882) );
  AND4X1_RVT U894 ( .A1(n884), .A2(n885), .A3(n886), .A4(n887), .Y(n816) );
  OR2X1_RVT U895 ( .A1(n888), .A2(n381), .Y(n887) );
  AND2X1_RVT U896 ( .A1(n889), .A2(n522), .Y(n888) );
  AND2X1_RVT U897 ( .A1(n890), .A2(n544), .Y(n889) );
  OR2X1_RVT U898 ( .A1(n156), .A2(n867), .Y(n544) );
  OR2X1_RVT U899 ( .A1(n12644), .A2(n478), .Y(n867) );
  OR2X1_RVT U900 ( .A1(n891), .A2(n12661), .Y(n886) );
  AND2X1_RVT U901 ( .A1(n892), .A2(n893), .Y(n891) );
  OR2X1_RVT U902 ( .A1(n894), .A2(n12803), .Y(n893) );
  AND2X1_RVT U903 ( .A1(n895), .A2(n896), .Y(n894) );
  OR2X1_RVT U904 ( .A1(n12643), .A2(n755), .Y(n896) );
  OR2X1_RVT U905 ( .A1(n12810), .A2(n401), .Y(n895) );
  AND2X1_RVT U906 ( .A1(n897), .A2(n898), .Y(n892) );
  OR2X1_RVT U907 ( .A1(n367), .A2(n899), .Y(n897) );
  OR2X1_RVT U908 ( .A1(n900), .A2(n401), .Y(n885) );
  AND4X1_RVT U909 ( .A1(n901), .A2(n902), .A3(n903), .A4(n367), .Y(n900) );
  OR2X1_RVT U910 ( .A1(n12811), .A2(n417), .Y(n903) );
  OR2X1_RVT U911 ( .A1(n12655), .A2(n436), .Y(n902) );
  OR2X1_RVT U912 ( .A1(n489), .A2(n467), .Y(n901) );
  OR2X1_RVT U913 ( .A1(n904), .A2(n343), .Y(n884) );
  AND4X1_RVT U914 ( .A1(n768), .A2(n905), .A3(n566), .A4(n482), .Y(n904) );
  OR2X1_RVT U915 ( .A1(n436), .A2(n899), .Y(n566) );
  OR2X1_RVT U916 ( .A1(n604), .A2(n811), .Y(n905) );
  OR2X1_RVT U917 ( .A1(n12649), .A2(n569), .Y(n768) );
  AND4X1_RVT U918 ( .A1(n907), .A2(n908), .A3(n909), .A4(n910), .Y(n906) );
  AND4X1_RVT U919 ( .A1(n419), .A2(n655), .A3(n911), .A4(n912), .Y(n910) );
  AND4X1_RVT U920 ( .A1(n734), .A2(n679), .A3(n824), .A4(n825), .Y(n912) );
  OR2X1_RVT U921 ( .A1(n827), .A2(n340), .Y(n825) );
  OR2X1_RVT U922 ( .A1(n12809), .A2(n458), .Y(n340) );
  OR2X1_RVT U923 ( .A1(n357), .A2(n866), .Y(n824) );
  OR2X1_RVT U924 ( .A1(n12814), .A2(n12663), .Y(n866) );
  OR2X1_RVT U925 ( .A1(n12803), .A2(n478), .Y(n357) );
  OR2X1_RVT U926 ( .A1(n12815), .A2(n376), .Y(n679) );
  OR2X1_RVT U927 ( .A1(n12672), .A2(n12656), .Y(n376) );
  OR2X1_RVT U928 ( .A1(n498), .A2(n913), .Y(n734) );
  OR2X1_RVT U929 ( .A1(n12663), .A2(n402), .Y(n913) );
  OR2X1_RVT U930 ( .A1(n400), .A2(n914), .Y(n911) );
  OR2X1_RVT U931 ( .A1(n528), .A2(n12654), .Y(n914) );
  OR2X1_RVT U932 ( .A1(n467), .A2(n915), .Y(n655) );
  OR2X1_RVT U933 ( .A1(n401), .A2(n12661), .Y(n915) );
  OR2X1_RVT U934 ( .A1(n12807), .A2(n826), .Y(n419) );
  OR2X1_RVT U935 ( .A1(n12656), .A2(n418), .Y(n826) );
  AND4X1_RVT U936 ( .A1(n916), .A2(n917), .A3(n918), .A4(n919), .Y(n909) );
  AND4X1_RVT U937 ( .A1(n920), .A2(n921), .A3(n922), .A4(n923), .Y(n919) );
  OR2X1_RVT U938 ( .A1(n434), .A2(n924), .Y(n923) );
  OR2X1_RVT U939 ( .A1(n12645), .A2(n504), .Y(n924) );
  OR2X1_RVT U940 ( .A1(n417), .A2(n925), .Y(n922) );
  OR2X1_RVT U941 ( .A1(n926), .A2(n381), .Y(n925) );
  AND2X1_RVT U942 ( .A1(n360), .A2(n420), .Y(n926) );
  OR2X1_RVT U943 ( .A1(n927), .A2(n928), .Y(n921) );
  AND2X1_RVT U944 ( .A1(n575), .A2(n531), .Y(n927) );
  OR2X1_RVT U945 ( .A1(n12808), .A2(n164), .Y(n531) );
  OR2X1_RVT U946 ( .A1(n12804), .A2(n12666), .Y(n575) );
  OR2X1_RVT U947 ( .A1(n929), .A2(n415), .Y(n920) );
  AND2X1_RVT U948 ( .A1(n811), .A2(n930), .Y(n929) );
  OR2X1_RVT U949 ( .A1(n12806), .A2(n156), .Y(n930) );
  OR2X1_RVT U950 ( .A1(n931), .A2(n12668), .Y(n918) );
  AND2X1_RVT U951 ( .A1(n802), .A2(n932), .Y(n931) );
  OR2X1_RVT U952 ( .A1(n408), .A2(n755), .Y(n932) );
  OR2X1_RVT U953 ( .A1(n12649), .A2(n620), .Y(n802) );
  OR2X1_RVT U954 ( .A1(n12810), .A2(n408), .Y(n620) );
  OR2X1_RVT U955 ( .A1(n933), .A2(n569), .Y(n917) );
  AND2X1_RVT U956 ( .A1(n522), .A2(n794), .Y(n933) );
  OR2X1_RVT U957 ( .A1(n378), .A2(n467), .Y(n522) );
  OR2X1_RVT U958 ( .A1(n934), .A2(n458), .Y(n916) );
  AND2X1_RVT U959 ( .A1(n421), .A2(n423), .Y(n934) );
  AND4X1_RVT U960 ( .A1(n935), .A2(n936), .A3(n937), .A4(n938), .Y(n908) );
  AND4X1_RVT U961 ( .A1(n939), .A2(n940), .A3(n941), .A4(n942), .Y(n938) );
  OR2X1_RVT U962 ( .A1(n943), .A2(n12652), .Y(n942) );
  AND2X1_RVT U963 ( .A1(n349), .A2(n641), .Y(n943) );
  OR2X1_RVT U964 ( .A1(n498), .A2(n529), .Y(n641) );
  OR2X1_RVT U965 ( .A1(n12655), .A2(n381), .Y(n529) );
  OR2X1_RVT U966 ( .A1(n12659), .A2(n944), .Y(n349) );
  OR2X1_RVT U967 ( .A1(n12642), .A2(n12648), .Y(n944) );
  OR2X1_RVT U968 ( .A1(n945), .A2(n12666), .Y(n941) );
  AND2X1_RVT U969 ( .A1(n658), .A2(n946), .Y(n945) );
  OR2X1_RVT U970 ( .A1(n12671), .A2(n154), .Y(n946) );
  OR2X1_RVT U971 ( .A1(n12669), .A2(n465), .Y(n658) );
  OR2X1_RVT U972 ( .A1(n947), .A2(n12647), .Y(n940) );
  AND2X1_RVT U973 ( .A1(n676), .A2(n948), .Y(n947) );
  OR2X1_RVT U974 ( .A1(n12672), .A2(n401), .Y(n948) );
  OR2X1_RVT U975 ( .A1(n343), .A2(n949), .Y(n676) );
  OR2X1_RVT U976 ( .A1(n950), .A2(n402), .Y(n939) );
  AND2X1_RVT U977 ( .A1(n951), .A2(n952), .Y(n950) );
  OR2X1_RVT U978 ( .A1(n458), .A2(n12669), .Y(n952) );
  AND2X1_RVT U979 ( .A1(n953), .A2(n434), .Y(n951) );
  OR2X1_RVT U980 ( .A1(n420), .A2(n381), .Y(n434) );
  OR2X1_RVT U981 ( .A1(n12644), .A2(n465), .Y(n953) );
  OR2X1_RVT U982 ( .A1(n12818), .A2(n420), .Y(n465) );
  OR2X1_RVT U983 ( .A1(n954), .A2(n478), .Y(n937) );
  AND4X1_RVT U984 ( .A1(n955), .A2(n956), .A3(n631), .A4(n541), .Y(n954) );
  OR2X1_RVT U985 ( .A1(n604), .A2(n704), .Y(n541) );
  OR2X1_RVT U986 ( .A1(n436), .A2(n883), .Y(n631) );
  OR2X1_RVT U987 ( .A1(n12650), .A2(n12643), .Y(n883) );
  OR2X1_RVT U988 ( .A1(n156), .A2(n358), .Y(n956) );
  OR2X1_RVT U989 ( .A1(n154), .A2(n12669), .Y(n955) );
  OR2X1_RVT U990 ( .A1(n957), .A2(n414), .Y(n936) );
  AND2X1_RVT U991 ( .A1(n958), .A2(n435), .Y(n957) );
  AND2X1_RVT U992 ( .A1(n890), .A2(n685), .Y(n958) );
  OR2X1_RVT U993 ( .A1(n959), .A2(n12815), .Y(n685) );
  AND2X1_RVT U994 ( .A1(n456), .A2(n960), .Y(n959) );
  OR2X1_RVT U995 ( .A1(n12647), .A2(n343), .Y(n960) );
  OR2X1_RVT U996 ( .A1(n504), .A2(n642), .Y(n890) );
  OR2X1_RVT U997 ( .A1(n489), .A2(n378), .Y(n642) );
  OR2X1_RVT U998 ( .A1(n961), .A2(n482), .Y(n935) );
  AND2X1_RVT U999 ( .A1(n962), .A2(n12655), .Y(n961) );
  AND2X1_RVT U1000 ( .A1(n963), .A2(n663), .Y(n962) );
  OR2X1_RVT U1001 ( .A1(n504), .A2(n604), .Y(n963) );
  AND4X1_RVT U1002 ( .A1(n964), .A2(n965), .A3(n966), .A4(n967), .Y(n907) );
  AND2X1_RVT U1003 ( .A1(n968), .A2(n969), .Y(n967) );
  OR2X1_RVT U1004 ( .A1(n12811), .A2(n584), .Y(n969) );
  OR2X1_RVT U1005 ( .A1(n12663), .A2(n970), .Y(n584) );
  OR2X1_RVT U1006 ( .A1(n400), .A2(n489), .Y(n970) );
  AND2X1_RVT U1007 ( .A1(n971), .A2(n972), .Y(n968) );
  OR2X1_RVT U1008 ( .A1(n373), .A2(n384), .Y(n972) );
  OR2X1_RVT U1009 ( .A1(n417), .A2(n612), .Y(n384) );
  OR2X1_RVT U1010 ( .A1(n12807), .A2(n378), .Y(n612) );
  OR2X1_RVT U1011 ( .A1(n420), .A2(n497), .Y(n971) );
  OR2X1_RVT U1012 ( .A1(n408), .A2(n973), .Y(n497) );
  OR2X1_RVT U1013 ( .A1(n408), .A2(n588), .Y(n966) );
  OR2X1_RVT U1014 ( .A1(n156), .A2(n12665), .Y(n588) );
  OR2X1_RVT U1015 ( .A1(n974), .A2(n364), .Y(n965) );
  AND4X1_RVT U1016 ( .A1(n975), .A2(n976), .A3(n977), .A4(n978), .Y(n974) );
  OR2X1_RVT U1017 ( .A1(n12805), .A2(n979), .Y(n977) );
  OR2X1_RVT U1018 ( .A1(n980), .A2(n12812), .Y(n979) );
  AND2X1_RVT U1019 ( .A1(n415), .A2(n981), .Y(n980) );
  OR2X1_RVT U1020 ( .A1(n12658), .A2(n982), .Y(n976) );
  OR2X1_RVT U1021 ( .A1(n721), .A2(n358), .Y(n982) );
  OR2X1_RVT U1022 ( .A1(n341), .A2(n367), .Y(n975) );
  OR2X1_RVT U1023 ( .A1(n12809), .A2(n467), .Y(n367) );
  OR2X1_RVT U1024 ( .A1(n841), .A2(n755), .Y(n964) );
  OR2X1_RVT U1025 ( .A1(n12674), .A2(n378), .Y(n755) );
  AND4X1_RVT U1026 ( .A1(n984), .A2(n985), .A3(n986), .A4(n987), .Y(n983) );
  AND4X1_RVT U1027 ( .A1(n988), .A2(n989), .A3(n990), .A4(n991), .Y(n987) );
  AND4X1_RVT U1028 ( .A1(n992), .A2(n993), .A3(n994), .A4(n995), .Y(n991) );
  OR2X1_RVT U1029 ( .A1(n829), .A2(n973), .Y(n995) );
  OR2X1_RVT U1030 ( .A1(n12808), .A2(n12668), .Y(n973) );
  OR2X1_RVT U1031 ( .A1(n12642), .A2(n12652), .Y(n829) );
  OR2X1_RVT U1032 ( .A1(n996), .A2(n415), .Y(n994) );
  AND2X1_RVT U1033 ( .A1(n361), .A2(n928), .Y(n996) );
  OR2X1_RVT U1034 ( .A1(n156), .A2(n997), .Y(n361) );
  OR2X1_RVT U1035 ( .A1(n12642), .A2(n12805), .Y(n997) );
  OR2X1_RVT U1036 ( .A1(n998), .A2(n343), .Y(n993) );
  OR2X1_RVT U1037 ( .A1(n12656), .A2(n504), .Y(n343) );
  AND2X1_RVT U1038 ( .A1(n479), .A2(n999), .Y(n998) );
  OR2X1_RVT U1039 ( .A1(n358), .A2(n560), .Y(n999) );
  OR2X1_RVT U1040 ( .A1(n12660), .A2(n12648), .Y(n358) );
  OR2X1_RVT U1041 ( .A1(n604), .A2(n1000), .Y(n479) );
  OR2X1_RVT U1042 ( .A1(n12816), .A2(n12663), .Y(n1000) );
  OR2X1_RVT U1043 ( .A1(n1001), .A2(n402), .Y(n992) );
  AND2X1_RVT U1044 ( .A1(n799), .A2(n1002), .Y(n1001) );
  OR2X1_RVT U1045 ( .A1(n1003), .A2(n12805), .Y(n1002) );
  AND2X1_RVT U1046 ( .A1(n458), .A2(n811), .Y(n1003) );
  OR2X1_RVT U1047 ( .A1(n12813), .A2(n420), .Y(n811) );
  OR2X1_RVT U1048 ( .A1(n12669), .A2(n1004), .Y(n799) );
  OR2X1_RVT U1049 ( .A1(n12818), .A2(n12814), .Y(n1004) );
  OR2X1_RVT U1050 ( .A1(n1005), .A2(n12647), .Y(n990) );
  AND2X1_RVT U1051 ( .A1(n1006), .A2(n1007), .Y(n1005) );
  OR2X1_RVT U1052 ( .A1(n1008), .A2(n504), .Y(n1007) );
  AND2X1_RVT U1053 ( .A1(n569), .A2(n1009), .Y(n1008) );
  OR2X1_RVT U1054 ( .A1(n360), .A2(n482), .Y(n1006) );
  OR2X1_RVT U1055 ( .A1(n12661), .A2(n418), .Y(n482) );
  OR2X1_RVT U1056 ( .A1(n1010), .A2(n12814), .Y(n989) );
  AND2X1_RVT U1057 ( .A1(n574), .A2(n733), .Y(n1010) );
  OR2X1_RVT U1058 ( .A1(n12659), .A2(n1011), .Y(n733) );
  OR2X1_RVT U1059 ( .A1(n414), .A2(n12648), .Y(n1011) );
  OR2X1_RVT U1060 ( .A1(n360), .A2(n841), .Y(n574) );
  OR2X1_RVT U1061 ( .A1(n12648), .A2(n12663), .Y(n841) );
  OR2X1_RVT U1062 ( .A1(n1012), .A2(n12645), .Y(n988) );
  AND2X1_RVT U1063 ( .A1(n614), .A2(n1013), .Y(n1012) );
  OR2X1_RVT U1064 ( .A1(n828), .A2(n408), .Y(n1013) );
  OR2X1_RVT U1065 ( .A1(n467), .A2(n949), .Y(n614) );
  OR2X1_RVT U1066 ( .A1(n12813), .A2(n156), .Y(n949) );
  AND2X1_RVT U1067 ( .A1(n12649), .A2(n12816), .Y(n710) );
  AND4X1_RVT U1068 ( .A1(n1014), .A2(n1015), .A3(n1016), .A4(n1017), .Y(n986)
         );
  AND4X1_RVT U1069 ( .A1(n1018), .A2(n1019), .A3(n1020), .A4(n1021), .Y(n1017)
         );
  OR2X1_RVT U1070 ( .A1(n1022), .A2(n12654), .Y(n1021) );
  AND2X1_RVT U1071 ( .A1(n601), .A2(n672), .Y(n1022) );
  OR2X1_RVT U1072 ( .A1(n417), .A2(n928), .Y(n672) );
  OR2X1_RVT U1073 ( .A1(n12816), .A2(n414), .Y(n928) );
  OR2X1_RVT U1074 ( .A1(n12803), .A2(n12644), .Y(n417) );
  OR2X1_RVT U1075 ( .A1(n12645), .A2(n704), .Y(n601) );
  OR2X1_RVT U1076 ( .A1(n12649), .A2(n12663), .Y(n704) );
  OR2X1_RVT U1077 ( .A1(n1023), .A2(n12812), .Y(n1020) );
  AND2X1_RVT U1078 ( .A1(n763), .A2(n1024), .Y(n1023) );
  OR2X1_RVT U1079 ( .A1(n721), .A2(n431), .Y(n1024) );
  OR2X1_RVT U1080 ( .A1(n604), .A2(n1025), .Y(n431) );
  OR2X1_RVT U1081 ( .A1(n12674), .A2(n12650), .Y(n1025) );
  OR2X1_RVT U1082 ( .A1(n12658), .A2(n1026), .Y(n763) );
  OR2X1_RVT U1083 ( .A1(n604), .A2(n400), .Y(n1026) );
  OR2X1_RVT U1084 ( .A1(n1027), .A2(n12818), .Y(n1019) );
  AND2X1_RVT U1085 ( .A1(n709), .A2(n638), .Y(n1027) );
  OR2X1_RVT U1086 ( .A1(n420), .A2(n456), .Y(n638) );
  OR2X1_RVT U1087 ( .A1(n12810), .A2(n604), .Y(n456) );
  OR2X1_RVT U1088 ( .A1(n828), .A2(n436), .Y(n709) );
  OR2X1_RVT U1089 ( .A1(n12655), .A2(n12815), .Y(n828) );
  OR2X1_RVT U1090 ( .A1(n1028), .A2(n478), .Y(n1018) );
  AND2X1_RVT U1091 ( .A1(n1029), .A2(n1030), .Y(n1028) );
  OR2X1_RVT U1092 ( .A1(n400), .A2(n827), .Y(n1030) );
  OR2X1_RVT U1093 ( .A1(n12812), .A2(n164), .Y(n827) );
  AND2X1_RVT U1094 ( .A1(n1031), .A2(n695), .Y(n1029) );
  OR2X1_RVT U1095 ( .A1(n408), .A2(n1032), .Y(n695) );
  OR2X1_RVT U1096 ( .A1(n12671), .A2(n12650), .Y(n1032) );
  OR2X1_RVT U1097 ( .A1(n464), .A2(n401), .Y(n1016) );
  OR2X1_RVT U1098 ( .A1(n12805), .A2(n360), .Y(n464) );
  OR2X1_RVT U1099 ( .A1(n1033), .A2(n364), .Y(n1015) );
  AND2X1_RVT U1100 ( .A1(n1034), .A2(n545), .Y(n1033) );
  AND2X1_RVT U1101 ( .A1(n1035), .A2(n1036), .Y(n545) );
  OR2X1_RVT U1102 ( .A1(n12659), .A2(n569), .Y(n1036) );
  OR2X1_RVT U1103 ( .A1(n467), .A2(n341), .Y(n1035) );
  OR2X1_RVT U1104 ( .A1(n12644), .A2(n414), .Y(n341) );
  AND2X1_RVT U1105 ( .A1(n1037), .A2(n731), .Y(n1034) );
  OR2X1_RVT U1106 ( .A1(n498), .A2(n981), .Y(n731) );
  OR2X1_RVT U1107 ( .A1(n12807), .A2(n154), .Y(n981) );
  OR2X1_RVT U1108 ( .A1(n360), .A2(n527), .Y(n1037) );
  OR2X1_RVT U1109 ( .A1(n12643), .A2(n1038), .Y(n527) );
  OR2X1_RVT U1110 ( .A1(n12803), .A2(n12672), .Y(n1038) );
  OR2X1_RVT U1111 ( .A1(n1039), .A2(n12803), .Y(n1014) );
  AND4X1_RVT U1112 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n873), .Y(n1039)
         );
  OR2X1_RVT U1113 ( .A1(n414), .A2(n794), .Y(n873) );
  OR2X1_RVT U1114 ( .A1(n12808), .A2(n12814), .Y(n794) );
  OR2X1_RVT U1115 ( .A1(n414), .A2(n1043), .Y(n1042) );
  OR2X1_RVT U1116 ( .A1(n12649), .A2(n12654), .Y(n1043) );
  OR2X1_RVT U1117 ( .A1(n12813), .A2(n373), .Y(n414) );
  OR2X1_RVT U1118 ( .A1(n1044), .A2(n495), .Y(n1041) );
  OR2X1_RVT U1119 ( .A1(n12643), .A2(n339), .Y(n495) );
  AND2X1_RVT U1120 ( .A1(n478), .A2(n1045), .Y(n1044) );
  OR2X1_RVT U1121 ( .A1(n12811), .A2(n378), .Y(n1045) );
  OR2X1_RVT U1122 ( .A1(n12807), .A2(n12654), .Y(n478) );
  OR2X1_RVT U1123 ( .A1(n12809), .A2(n1009), .Y(n1040) );
  OR2X1_RVT U1124 ( .A1(n12813), .A2(n418), .Y(n1009) );
  OR2X1_RVT U1125 ( .A1(n364), .A2(n154), .Y(n418) );
  AND4X1_RVT U1126 ( .A1(n1046), .A2(n1047), .A3(n1048), .A4(n1049), .Y(n985)
         );
  AND4X1_RVT U1127 ( .A1(n1050), .A2(n1051), .A3(n1052), .A4(n1053), .Y(n1049)
         );
  OR2X1_RVT U1128 ( .A1(n436), .A2(n563), .Y(n1053) );
  OR2X1_RVT U1129 ( .A1(n12656), .A2(n458), .Y(n563) );
  OR2X1_RVT U1130 ( .A1(n12660), .A2(n604), .Y(n436) );
  OR2X1_RVT U1131 ( .A1(n423), .A2(n899), .Y(n1052) );
  OR2X1_RVT U1132 ( .A1(n12817), .A2(n12643), .Y(n899) );
  OR2X1_RVT U1133 ( .A1(n489), .A2(n415), .Y(n423) );
  OR2X1_RVT U1134 ( .A1(n408), .A2(n435), .Y(n1051) );
  OR2X1_RVT U1135 ( .A1(n12652), .A2(n12665), .Y(n435) );
  OR2X1_RVT U1136 ( .A1(n12642), .A2(n12804), .Y(n408) );
  OR2X1_RVT U1137 ( .A1(n164), .A2(n774), .Y(n1050) );
  OR2X1_RVT U1138 ( .A1(n12650), .A2(n561), .Y(n774) );
  OR2X1_RVT U1139 ( .A1(n378), .A2(n808), .Y(n1048) );
  OR2X1_RVT U1140 ( .A1(n164), .A2(n1054), .Y(n808) );
  OR2X1_RVT U1141 ( .A1(n12810), .A2(n12663), .Y(n1054) );
  AND2X1_RVT U1142 ( .A1(n12644), .A2(n12647), .Y(n838) );
  OR2X1_RVT U1143 ( .A1(n420), .A2(n368), .Y(n1047) );
  OR2X1_RVT U1144 ( .A1(n12672), .A2(n1055), .Y(n368) );
  OR2X1_RVT U1145 ( .A1(n12811), .A2(n12803), .Y(n1055) );
  OR2X1_RVT U1146 ( .A1(n12649), .A2(n400), .Y(n420) );
  OR2X1_RVT U1147 ( .A1(n467), .A2(n1031), .Y(n1046) );
  OR2X1_RVT U1148 ( .A1(n12645), .A2(n422), .Y(n1031) );
  OR2X1_RVT U1149 ( .A1(n12813), .A2(n12814), .Y(n422) );
  AND4X1_RVT U1150 ( .A1(n1056), .A2(n533), .A3(n1057), .A4(n1058), .Y(n984)
         );
  OR2X1_RVT U1151 ( .A1(n12649), .A2(n978), .Y(n1058) );
  OR2X1_RVT U1152 ( .A1(n12809), .A2(n528), .Y(n978) );
  OR2X1_RVT U1153 ( .A1(n12647), .A2(n569), .Y(n528) );
  OR2X1_RVT U1154 ( .A1(n12642), .A2(n395), .Y(n569) );
  AND2X1_RVT U1155 ( .A1(n1059), .A2(n1060), .Y(n1057) );
  OR2X1_RVT U1156 ( .A1(n12671), .A2(n898), .Y(n1060) );
  OR2X1_RVT U1157 ( .A1(n467), .A2(n560), .Y(n898) );
  OR2X1_RVT U1158 ( .A1(n12649), .A2(n12643), .Y(n560) );
  OR2X1_RVT U1159 ( .A1(n12644), .A2(n356), .Y(n395) );
  OR2X1_RVT U1160 ( .A1(n12816), .A2(n629), .Y(n1059) );
  OR2X1_RVT U1161 ( .A1(n12668), .A2(n663), .Y(n629) );
  OR2X1_RVT U1162 ( .A1(n12808), .A2(n12803), .Y(n663) );
  OR2X1_RVT U1163 ( .A1(n12806), .A2(n12660), .Y(n339) );
  AND2X1_RVT U1164 ( .A1(n1061), .A2(n1062), .Y(n533) );
  OR2X1_RVT U1165 ( .A1(n415), .A2(n401), .Y(n1062) );
  OR2X1_RVT U1166 ( .A1(n12815), .A2(n373), .Y(n401) );
  AND2X1_RVT U1167 ( .A1(n400), .A2(n364), .Y(n453) );
  OR2X1_RVT U1168 ( .A1(n12655), .A2(n467), .Y(n415) );
  OR2X1_RVT U1169 ( .A1(n12804), .A2(n504), .Y(n467) );
  OR2X1_RVT U1170 ( .A1(n1063), .A2(n458), .Y(n1061) );
  OR2X1_RVT U1171 ( .A1(n12649), .A2(n154), .Y(n458) );
  AND2X1_RVT U1172 ( .A1(n12817), .A2(n12642), .Y(n721) );
  OR2X1_RVT U1173 ( .A1(n12648), .A2(n561), .Y(n1063) );
  OR2X1_RVT U1174 ( .A1(n12813), .A2(n12665), .Y(n561) );
  AND2X1_RVT U1175 ( .A1(n1064), .A2(n1065), .Y(n1056) );
  OR2X1_RVT U1176 ( .A1(n381), .A2(n714), .Y(n1065) );
  OR2X1_RVT U1177 ( .A1(n12650), .A2(n421), .Y(n714) );
  OR2X1_RVT U1178 ( .A1(n12665), .A2(n498), .Y(n421) );
  OR2X1_RVT U1179 ( .A1(n12645), .A2(n12648), .Y(n498) );
  OR2X1_RVT U1180 ( .A1(n12810), .A2(n12808), .Y(n360) );
  OR2X1_RVT U1181 ( .A1(n12818), .A2(n12812), .Y(n381) );
  XOR2X1_RVT U1182 ( .A1(key[68]), .A2(state[68]), .Y(n356) );
  OR2X1_RVT U1183 ( .A1(n373), .A2(n502), .Y(n1064) );
  OR2X1_RVT U1184 ( .A1(n604), .A2(n795), .Y(n502) );
  OR2X1_RVT U1185 ( .A1(n12652), .A2(n402), .Y(n795) );
  OR2X1_RVT U1186 ( .A1(n12811), .A2(n504), .Y(n402) );
  XOR2X1_RVT U1187 ( .A1(key[66]), .A2(state[66]), .Y(n504) );
  XOR2X1_RVT U1188 ( .A1(key[67]), .A2(state[67]), .Y(n438) );
  OR2X1_RVT U1189 ( .A1(n12816), .A2(n12650), .Y(n378) );
  XOR2X1_RVT U1190 ( .A1(key[69]), .A2(state[69]), .Y(n364) );
  XOR2X1_RVT U1191 ( .A1(key[70]), .A2(state[70]), .Y(n400) );
  OR2X1_RVT U1192 ( .A1(n12806), .A2(n12648), .Y(n604) );
  XOR2X1_RVT U1193 ( .A1(key[64]), .A2(state[64]), .Y(n379) );
  XOR2X1_RVT U1194 ( .A1(key[65]), .A2(state[65]), .Y(n489) );
  XOR2X1_RVT U1195 ( .A1(key[71]), .A2(state[71]), .Y(n373) );
  AND4X1_RVT U1196 ( .A1(n1067), .A2(n1068), .A3(n1069), .A4(n1070), .Y(n1066)
         );
  AND4X1_RVT U1197 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .Y(n1070)
         );
  AND4X1_RVT U1198 ( .A1(n1075), .A2(n1076), .A3(n1077), .A4(n1078), .Y(n1074)
         );
  OR2X1_RVT U1199 ( .A1(n12636), .A2(n1080), .Y(n1073) );
  OR2X1_RVT U1200 ( .A1(n1081), .A2(n1082), .Y(n1071) );
  OR2X1_RVT U1201 ( .A1(n12923), .A2(n1083), .Y(n1082) );
  AND4X1_RVT U1202 ( .A1(n1084), .A2(n1085), .A3(n1086), .A4(n1087), .Y(n1069)
         );
  OR2X1_RVT U1203 ( .A1(n1088), .A2(n12921), .Y(n1087) );
  AND2X1_RVT U1204 ( .A1(n1089), .A2(n1090), .Y(n1088) );
  AND2X1_RVT U1205 ( .A1(n1091), .A2(n1092), .Y(n1086) );
  OR2X1_RVT U1206 ( .A1(n1093), .A2(n11), .Y(n1092) );
  AND2X1_RVT U1207 ( .A1(n1094), .A2(n1095), .Y(n1093) );
  OR2X1_RVT U1208 ( .A1(n12627), .A2(n1097), .Y(n1095) );
  OR2X1_RVT U1209 ( .A1(n1083), .A2(n1098), .Y(n1094) );
  OR2X1_RVT U1210 ( .A1(n1099), .A2(n12633), .Y(n1091) );
  AND2X1_RVT U1211 ( .A1(n1101), .A2(n1102), .Y(n1099) );
  OR2X1_RVT U1212 ( .A1(n1103), .A2(n1104), .Y(n1085) );
  AND2X1_RVT U1213 ( .A1(n1105), .A2(n1106), .Y(n1103) );
  OR2X1_RVT U1214 ( .A1(n12628), .A2(n1107), .Y(n1106) );
  AND2X1_RVT U1215 ( .A1(n1108), .A2(n1109), .Y(n1105) );
  AND2X1_RVT U1216 ( .A1(n1110), .A2(n1111), .Y(n1084) );
  OR2X1_RVT U1217 ( .A1(n1112), .A2(n12610), .Y(n1111) );
  AND2X1_RVT U1218 ( .A1(n1114), .A2(n1115), .Y(n1112) );
  OR2X1_RVT U1219 ( .A1(n1116), .A2(n1117), .Y(n1115) );
  OR2X1_RVT U1220 ( .A1(n12619), .A2(n12614), .Y(n1117) );
  OR2X1_RVT U1221 ( .A1(n1120), .A2(n1121), .Y(n1110) );
  AND2X1_RVT U1222 ( .A1(n1122), .A2(n1123), .Y(n1120) );
  AND2X1_RVT U1223 ( .A1(n1124), .A2(n1125), .Y(n1122) );
  AND4X1_RVT U1224 ( .A1(n1126), .A2(n1127), .A3(n1128), .A4(n1129), .Y(n1068)
         );
  AND4X1_RVT U1225 ( .A1(n1130), .A2(n1131), .A3(n1132), .A4(n1133), .Y(n1129)
         );
  OR2X1_RVT U1226 ( .A1(n1134), .A2(n12639), .Y(n1133) );
  AND4X1_RVT U1227 ( .A1(n1136), .A2(n1137), .A3(n1138), .A4(n1139), .Y(n1134)
         );
  OR2X1_RVT U1228 ( .A1(n1140), .A2(n1107), .Y(n1139) );
  OR2X1_RVT U1229 ( .A1(n1141), .A2(n12625), .Y(n1138) );
  OR2X1_RVT U1230 ( .A1(n1143), .A2(n12616), .Y(n1132) );
  AND4X1_RVT U1231 ( .A1(n1144), .A2(n1145), .A3(n1146), .A4(n1147), .Y(n1143)
         );
  OR2X1_RVT U1232 ( .A1(n1148), .A2(n1149), .Y(n1147) );
  OR2X1_RVT U1233 ( .A1(n12633), .A2(n12628), .Y(n1149) );
  AND2X1_RVT U1234 ( .A1(n1150), .A2(n1151), .Y(n1146) );
  OR2X1_RVT U1235 ( .A1(n12925), .A2(n1152), .Y(n1145) );
  OR2X1_RVT U1236 ( .A1(n1153), .A2(n1154), .Y(n1144) );
  AND2X1_RVT U1237 ( .A1(n1155), .A2(n1156), .Y(n1153) );
  OR2X1_RVT U1238 ( .A1(n12633), .A2(n1157), .Y(n1156) );
  OR2X1_RVT U1239 ( .A1(n1090), .A2(n1158), .Y(n1131) );
  OR2X1_RVT U1240 ( .A1(n1157), .A2(n1159), .Y(n1130) );
  OR2X1_RVT U1241 ( .A1(n1160), .A2(n1161), .Y(n1128) );
  OR2X1_RVT U1242 ( .A1(n1162), .A2(n1155), .Y(n1127) );
  OR2X1_RVT U1243 ( .A1(n1163), .A2(n1164), .Y(n1126) );
  AND4X1_RVT U1244 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .Y(n1067)
         );
  AND2X1_RVT U1245 ( .A1(n1169), .A2(n1170), .Y(n1168) );
  OR2X1_RVT U1246 ( .A1(n1154), .A2(n1171), .Y(n1170) );
  AND2X1_RVT U1247 ( .A1(n1172), .A2(n1173), .Y(n1169) );
  OR2X1_RVT U1248 ( .A1(n1174), .A2(n1097), .Y(n1173) );
  OR2X1_RVT U1249 ( .A1(n1098), .A2(n1175), .Y(n1172) );
  OR2X1_RVT U1250 ( .A1(n9), .A2(n1176), .Y(n1167) );
  OR2X1_RVT U1251 ( .A1(n1177), .A2(n12623), .Y(n1166) );
  OR2X1_RVT U1252 ( .A1(n12626), .A2(n1179), .Y(n1165) );
  AND4X1_RVT U1253 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .Y(n1180)
         );
  AND4X1_RVT U1254 ( .A1(n1185), .A2(n1076), .A3(n1186), .A4(n1187), .Y(n1184)
         );
  AND4X1_RVT U1255 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .Y(n1187)
         );
  OR2X1_RVT U1256 ( .A1(n1097), .A2(n1192), .Y(n1191) );
  OR2X1_RVT U1257 ( .A1(n1193), .A2(n12638), .Y(n1192) );
  OR2X1_RVT U1258 ( .A1(n1098), .A2(n1194), .Y(n1190) );
  OR2X1_RVT U1259 ( .A1(n9), .A2(n12622), .Y(n1194) );
  OR2X1_RVT U1260 ( .A1(n1195), .A2(n1141), .Y(n1189) );
  AND2X1_RVT U1261 ( .A1(n1152), .A2(n1196), .Y(n1195) );
  OR2X1_RVT U1262 ( .A1(n1197), .A2(n1198), .Y(n1188) );
  AND2X1_RVT U1263 ( .A1(n1199), .A2(n1200), .Y(n1197) );
  AND2X1_RVT U1264 ( .A1(n1201), .A2(n1202), .Y(n1186) );
  OR2X1_RVT U1265 ( .A1(n1148), .A2(n1203), .Y(n1202) );
  OR2X1_RVT U1266 ( .A1(n1204), .A2(n12923), .Y(n1203) );
  OR2X1_RVT U1267 ( .A1(n1205), .A2(n1206), .Y(n1201) );
  OR2X1_RVT U1268 ( .A1(n1207), .A2(n12627), .Y(n1206) );
  OR2X1_RVT U1269 ( .A1(n1083), .A2(n1208), .Y(n1076) );
  AND4X1_RVT U1270 ( .A1(n1209), .A2(n1210), .A3(n1211), .A4(n1212), .Y(n1183)
         );
  AND4X1_RVT U1271 ( .A1(n1213), .A2(n1214), .A3(n1215), .A4(n1216), .Y(n1212)
         );
  OR2X1_RVT U1272 ( .A1(n1217), .A2(n12641), .Y(n1216) );
  AND2X1_RVT U1273 ( .A1(n1219), .A2(n1220), .Y(n1217) );
  OR2X1_RVT U1274 ( .A1(n12610), .A2(n1098), .Y(n1220) );
  OR2X1_RVT U1275 ( .A1(n1221), .A2(n1100), .Y(n1215) );
  AND2X1_RVT U1276 ( .A1(n1222), .A2(n1223), .Y(n1221) );
  OR2X1_RVT U1277 ( .A1(n1224), .A2(n12922), .Y(n1214) );
  AND2X1_RVT U1278 ( .A1(n1225), .A2(n1226), .Y(n1224) );
  OR2X1_RVT U1279 ( .A1(n1227), .A2(n1176), .Y(n1226) );
  AND2X1_RVT U1280 ( .A1(n12641), .A2(n12625), .Y(n1227) );
  OR2X1_RVT U1281 ( .A1(n1228), .A2(n12611), .Y(n1213) );
  AND2X1_RVT U1282 ( .A1(n1230), .A2(n1231), .Y(n1228) );
  OR2X1_RVT U1283 ( .A1(n1232), .A2(n12617), .Y(n1211) );
  AND2X1_RVT U1284 ( .A1(n1233), .A2(n1234), .Y(n1232) );
  OR2X1_RVT U1285 ( .A1(n12625), .A2(n1235), .Y(n1234) );
  AND2X1_RVT U1286 ( .A1(n1236), .A2(n1237), .Y(n1233) );
  OR2X1_RVT U1287 ( .A1(n1238), .A2(n1239), .Y(n1236) );
  OR2X1_RVT U1288 ( .A1(n1083), .A2(n1154), .Y(n1239) );
  OR2X1_RVT U1289 ( .A1(n1240), .A2(n12919), .Y(n1210) );
  AND2X1_RVT U1290 ( .A1(n1241), .A2(n1242), .Y(n1240) );
  OR2X1_RVT U1291 ( .A1(n1243), .A2(n1244), .Y(n1209) );
  AND2X1_RVT U1292 ( .A1(n1245), .A2(n1246), .Y(n1243) );
  AND2X1_RVT U1293 ( .A1(n1247), .A2(n1248), .Y(n1245) );
  OR2X1_RVT U1294 ( .A1(n11), .A2(n1176), .Y(n1248) );
  OR2X1_RVT U1295 ( .A1(n12635), .A2(n1141), .Y(n1247) );
  AND4X1_RVT U1296 ( .A1(n1249), .A2(n1250), .A3(n1251), .A4(n1252), .Y(n1182)
         );
  AND4X1_RVT U1297 ( .A1(n1253), .A2(n1254), .A3(n1255), .A4(n1256), .Y(n1252)
         );
  OR2X1_RVT U1298 ( .A1(n1176), .A2(n1175), .Y(n1256) );
  OR2X1_RVT U1299 ( .A1(n1107), .A2(n1257), .Y(n1255) );
  OR2X1_RVT U1300 ( .A1(n1140), .A2(n1258), .Y(n1254) );
  OR2X1_RVT U1301 ( .A1(n1083), .A2(n1259), .Y(n1253) );
  AND2X1_RVT U1302 ( .A1(n1260), .A2(n1261), .Y(n1251) );
  OR2X1_RVT U1303 ( .A1(n12636), .A2(n1262), .Y(n1261) );
  OR2X1_RVT U1304 ( .A1(n12615), .A2(n1159), .Y(n1260) );
  OR2X1_RVT U1305 ( .A1(n1263), .A2(n1118), .Y(n1250) );
  AND4X1_RVT U1306 ( .A1(n1264), .A2(n1265), .A3(n1266), .A4(n1267), .Y(n1263)
         );
  OR2X1_RVT U1307 ( .A1(n1268), .A2(n1083), .Y(n1266) );
  OR2X1_RVT U1308 ( .A1(n12911), .A2(n1269), .Y(n1265) );
  OR2X1_RVT U1309 ( .A1(n1270), .A2(n12919), .Y(n1264) );
  AND2X1_RVT U1310 ( .A1(n1161), .A2(n1271), .Y(n1270) );
  OR2X1_RVT U1311 ( .A1(n1163), .A2(n1272), .Y(n1249) );
  AND4X1_RVT U1312 ( .A1(n1273), .A2(n1274), .A3(n1275), .A4(n1276), .Y(n1181)
         );
  AND4X1_RVT U1313 ( .A1(n1277), .A2(n1278), .A3(n1279), .A4(n1280), .Y(n1276)
         );
  OR2X1_RVT U1314 ( .A1(n12915), .A2(n1281), .Y(n1280) );
  OR2X1_RVT U1315 ( .A1(n12916), .A2(n1282), .Y(n1279) );
  OR2X1_RVT U1316 ( .A1(n12913), .A2(n1283), .Y(n1278) );
  OR2X1_RVT U1317 ( .A1(n12609), .A2(n1284), .Y(n1277) );
  OR2X1_RVT U1318 ( .A1(n1285), .A2(n12616), .Y(n1274) );
  AND4X1_RVT U1319 ( .A1(n1287), .A2(n1288), .A3(n1289), .A4(n1290), .Y(n1286)
         );
  AND4X1_RVT U1320 ( .A1(n1291), .A2(n1292), .A3(n1293), .A4(n1294), .Y(n1290)
         );
  AND4X1_RVT U1321 ( .A1(n1295), .A2(n1296), .A3(n1297), .A4(n1298), .Y(n1294)
         );
  OR2X1_RVT U1322 ( .A1(n1299), .A2(n12204), .Y(n1297) );
  AND2X1_RVT U1323 ( .A1(n1301), .A2(n1302), .Y(n1299) );
  OR2X1_RVT U1324 ( .A1(n1303), .A2(n12184), .Y(n1296) );
  AND2X1_RVT U1325 ( .A1(n1304), .A2(n1305), .Y(n1303) );
  OR2X1_RVT U1326 ( .A1(n1306), .A2(n12201), .Y(n1305) );
  OR2X1_RVT U1327 ( .A1(n1308), .A2(n12189), .Y(n1295) );
  AND2X1_RVT U1328 ( .A1(n1310), .A2(n1311), .Y(n1308) );
  OR2X1_RVT U1329 ( .A1(n1312), .A2(n1313), .Y(n1311) );
  OR2X1_RVT U1330 ( .A1(n1306), .A2(n12926), .Y(n1310) );
  OR2X1_RVT U1331 ( .A1(n1315), .A2(n85), .Y(n1293) );
  AND2X1_RVT U1332 ( .A1(n1316), .A2(n1317), .Y(n1315) );
  AND2X1_RVT U1333 ( .A1(n1318), .A2(n1319), .Y(n1316) );
  OR2X1_RVT U1334 ( .A1(n1320), .A2(n12871), .Y(n1292) );
  AND2X1_RVT U1335 ( .A1(n1321), .A2(n1322), .Y(n1320) );
  OR2X1_RVT U1336 ( .A1(n83), .A2(n1323), .Y(n1322) );
  OR2X1_RVT U1337 ( .A1(n1324), .A2(n1325), .Y(n1291) );
  AND2X1_RVT U1338 ( .A1(n1326), .A2(n1327), .Y(n1324) );
  OR2X1_RVT U1339 ( .A1(n1328), .A2(n1329), .Y(n1327) );
  AND2X1_RVT U1340 ( .A1(n1330), .A2(n1331), .Y(n1326) );
  OR2X1_RVT U1341 ( .A1(n1332), .A2(n1333), .Y(n1330) );
  OR2X1_RVT U1342 ( .A1(n12873), .A2(n1334), .Y(n1333) );
  AND4X1_RVT U1343 ( .A1(n1335), .A2(n1336), .A3(n1337), .A4(n1338), .Y(n1289)
         );
  AND2X1_RVT U1344 ( .A1(n1339), .A2(n1340), .Y(n1338) );
  OR2X1_RVT U1345 ( .A1(n1341), .A2(n1342), .Y(n1340) );
  AND2X1_RVT U1346 ( .A1(n1343), .A2(n1344), .Y(n1339) );
  OR2X1_RVT U1347 ( .A1(n1345), .A2(n1346), .Y(n1344) );
  OR2X1_RVT U1348 ( .A1(n1347), .A2(n1348), .Y(n1343) );
  OR2X1_RVT U1349 ( .A1(n1349), .A2(n1350), .Y(n1337) );
  AND4X1_RVT U1350 ( .A1(n1351), .A2(n1352), .A3(n1353), .A4(n1354), .Y(n1349)
         );
  OR2X1_RVT U1351 ( .A1(n12926), .A2(n1355), .Y(n1354) );
  OR2X1_RVT U1352 ( .A1(n12212), .A2(n83), .Y(n1355) );
  AND2X1_RVT U1353 ( .A1(n1357), .A2(n1358), .Y(n1353) );
  OR2X1_RVT U1354 ( .A1(n1359), .A2(n1360), .Y(n1357) );
  OR2X1_RVT U1355 ( .A1(n1361), .A2(n12150), .Y(n1360) );
  OR2X1_RVT U1356 ( .A1(n12871), .A2(n1313), .Y(n1352) );
  OR2X1_RVT U1357 ( .A1(n1362), .A2(n12150), .Y(n1336) );
  AND2X1_RVT U1358 ( .A1(n1363), .A2(n1364), .Y(n1362) );
  OR2X1_RVT U1359 ( .A1(n1365), .A2(n1332), .Y(n1364) );
  AND2X1_RVT U1360 ( .A1(n1366), .A2(n1367), .Y(n1363) );
  OR2X1_RVT U1361 ( .A1(n1368), .A2(n12875), .Y(n1335) );
  AND4X1_RVT U1362 ( .A1(n1369), .A2(n1370), .A3(n1371), .A4(n1372), .Y(n1368)
         );
  AND2X1_RVT U1363 ( .A1(n1373), .A2(n1374), .Y(n1371) );
  OR2X1_RVT U1364 ( .A1(n12186), .A2(n1376), .Y(n1369) );
  AND4X1_RVT U1365 ( .A1(n1377), .A2(n1378), .A3(n1379), .A4(n1380), .Y(n1288)
         );
  AND4X1_RVT U1366 ( .A1(n1381), .A2(n1382), .A3(n1383), .A4(n1384), .Y(n1380)
         );
  OR2X1_RVT U1367 ( .A1(n1332), .A2(n1385), .Y(n1384) );
  OR2X1_RVT U1368 ( .A1(n1386), .A2(n1387), .Y(n1383) );
  OR2X1_RVT U1369 ( .A1(n73), .A2(n1331), .Y(n1382) );
  OR2X1_RVT U1370 ( .A1(n72), .A2(n1370), .Y(n1381) );
  OR2X1_RVT U1371 ( .A1(n12206), .A2(n1389), .Y(n1379) );
  OR2X1_RVT U1372 ( .A1(n1314), .A2(n1390), .Y(n1378) );
  OR2X1_RVT U1373 ( .A1(n1391), .A2(n1392), .Y(n1377) );
  AND4X1_RVT U1374 ( .A1(n1393), .A2(n1394), .A3(n1395), .A4(n1396), .Y(n1287)
         );
  OR2X1_RVT U1375 ( .A1(n12870), .A2(n1397), .Y(n1396) );
  AND2X1_RVT U1376 ( .A1(n1398), .A2(n1399), .Y(n1395) );
  OR2X1_RVT U1377 ( .A1(n1356), .A2(n1400), .Y(n1399) );
  OR2X1_RVT U1378 ( .A1(n12874), .A2(n1401), .Y(n1398) );
  AND2X1_RVT U1379 ( .A1(n1402), .A2(n1403), .Y(n1393) );
  OR2X1_RVT U1380 ( .A1(n12868), .A2(n1404), .Y(n1403) );
  OR2X1_RVT U1381 ( .A1(n1307), .A2(n1301), .Y(n1402) );
  AND4X1_RVT U1382 ( .A1(n1406), .A2(n1407), .A3(n1408), .A4(n1409), .Y(n1405)
         );
  AND4X1_RVT U1383 ( .A1(n1410), .A2(n1411), .A3(n1412), .A4(n1413), .Y(n1409)
         );
  AND4X1_RVT U1384 ( .A1(n1414), .A2(n1072), .A3(n1242), .A4(n1415), .Y(n1413)
         );
  OR2X1_RVT U1385 ( .A1(n1416), .A2(n12910), .Y(n1072) );
  AND2X1_RVT U1386 ( .A1(n1417), .A2(n1418), .Y(n1416) );
  OR2X1_RVT U1387 ( .A1(n1116), .A2(n1419), .Y(n1418) );
  OR2X1_RVT U1388 ( .A1(n1420), .A2(n1198), .Y(n1417) );
  OR2X1_RVT U1389 ( .A1(n1421), .A2(n1157), .Y(n1414) );
  AND2X1_RVT U1390 ( .A1(n1422), .A2(n1423), .Y(n1421) );
  OR2X1_RVT U1391 ( .A1(n12915), .A2(n1141), .Y(n1423) );
  OR2X1_RVT U1392 ( .A1(n1424), .A2(n1100), .Y(n1412) );
  AND2X1_RVT U1393 ( .A1(n1425), .A2(n1426), .Y(n1424) );
  OR2X1_RVT U1394 ( .A1(n1427), .A2(n12921), .Y(n1426) );
  AND2X1_RVT U1395 ( .A1(n1148), .A2(n1428), .Y(n1427) );
  OR2X1_RVT U1396 ( .A1(n1429), .A2(n12636), .Y(n1411) );
  AND2X1_RVT U1397 ( .A1(n1430), .A2(n1431), .Y(n1429) );
  OR2X1_RVT U1398 ( .A1(n1141), .A2(n1107), .Y(n1431) );
  OR2X1_RVT U1399 ( .A1(n1432), .A2(n12619), .Y(n1410) );
  AND2X1_RVT U1400 ( .A1(n1225), .A2(n1433), .Y(n1432) );
  OR2X1_RVT U1401 ( .A1(n1154), .A2(n1434), .Y(n1225) );
  AND4X1_RVT U1402 ( .A1(n1435), .A2(n1436), .A3(n1437), .A4(n1438), .Y(n1408)
         );
  OR2X1_RVT U1403 ( .A1(n1439), .A2(n12626), .Y(n1438) );
  AND2X1_RVT U1404 ( .A1(n1440), .A2(n1441), .Y(n1439) );
  OR2X1_RVT U1405 ( .A1(n1198), .A2(n1098), .Y(n1441) );
  AND2X1_RVT U1406 ( .A1(n1442), .A2(n1443), .Y(n1440) );
  OR2X1_RVT U1407 ( .A1(n1238), .A2(n1419), .Y(n1442) );
  AND2X1_RVT U1408 ( .A1(n1444), .A2(n1445), .Y(n1437) );
  OR2X1_RVT U1409 ( .A1(n1446), .A2(n1229), .Y(n1445) );
  AND2X1_RVT U1410 ( .A1(n1447), .A2(n1137), .Y(n1446) );
  OR2X1_RVT U1411 ( .A1(n1083), .A2(n1198), .Y(n1137) );
  OR2X1_RVT U1412 ( .A1(n1448), .A2(n11), .Y(n1444) );
  AND2X1_RVT U1413 ( .A1(n1449), .A2(n1450), .Y(n1448) );
  OR2X1_RVT U1414 ( .A1(n1451), .A2(n12628), .Y(n1450) );
  AND2X1_RVT U1415 ( .A1(n1452), .A2(n1453), .Y(n1451) );
  OR2X1_RVT U1416 ( .A1(n12623), .A2(n1148), .Y(n1453) );
  OR2X1_RVT U1417 ( .A1(n12925), .A2(n12625), .Y(n1452) );
  AND2X1_RVT U1418 ( .A1(n1199), .A2(n1428), .Y(n1449) );
  OR2X1_RVT U1419 ( .A1(n1229), .A2(n1454), .Y(n1199) );
  OR2X1_RVT U1420 ( .A1(n12920), .A2(n12916), .Y(n1454) );
  OR2X1_RVT U1421 ( .A1(n1455), .A2(n1218), .Y(n1436) );
  AND4X1_RVT U1422 ( .A1(n1177), .A2(n1456), .A3(n1457), .A4(n1458), .Y(n1455)
         );
  OR2X1_RVT U1423 ( .A1(n12627), .A2(n1198), .Y(n1458) );
  AND2X1_RVT U1424 ( .A1(n1459), .A2(n1460), .Y(n1457) );
  OR2X1_RVT U1425 ( .A1(n12925), .A2(n12636), .Y(n1456) );
  AND2X1_RVT U1426 ( .A1(n1461), .A2(n1462), .Y(n1177) );
  OR2X1_RVT U1427 ( .A1(n1463), .A2(n9), .Y(n1462) );
  OR2X1_RVT U1428 ( .A1(n1141), .A2(n12910), .Y(n1461) );
  AND2X1_RVT U1429 ( .A1(n1464), .A2(n1465), .Y(n1435) );
  OR2X1_RVT U1430 ( .A1(n1466), .A2(n12912), .Y(n1465) );
  AND2X1_RVT U1431 ( .A1(n1467), .A2(n1468), .Y(n1466) );
  OR2X1_RVT U1432 ( .A1(n1469), .A2(n12630), .Y(n1468) );
  AND2X1_RVT U1433 ( .A1(n1470), .A2(n1471), .Y(n1469) );
  AND2X1_RVT U1434 ( .A1(n1472), .A2(n1473), .Y(n1467) );
  OR2X1_RVT U1435 ( .A1(n1474), .A2(n12639), .Y(n1464) );
  AND4X1_RVT U1436 ( .A1(n1475), .A2(n1476), .A3(n1477), .A4(n1478), .Y(n1474)
         );
  OR2X1_RVT U1437 ( .A1(n12924), .A2(n1479), .Y(n1477) );
  OR2X1_RVT U1438 ( .A1(n9), .A2(n1155), .Y(n1476) );
  OR2X1_RVT U1439 ( .A1(n1244), .A2(n1198), .Y(n1475) );
  AND4X1_RVT U1440 ( .A1(n1480), .A2(n1481), .A3(n1482), .A4(n1483), .Y(n1407)
         );
  AND2X1_RVT U1441 ( .A1(n1484), .A2(n1208), .Y(n1483) );
  OR2X1_RVT U1442 ( .A1(n12614), .A2(n1174), .Y(n1208) );
  AND2X1_RVT U1443 ( .A1(n1485), .A2(n1486), .Y(n1484) );
  OR2X1_RVT U1444 ( .A1(n1487), .A2(n1123), .Y(n1486) );
  OR2X1_RVT U1445 ( .A1(n1175), .A2(n1235), .Y(n1485) );
  OR2X1_RVT U1446 ( .A1(n9), .A2(n1488), .Y(n1482) );
  OR2X1_RVT U1447 ( .A1(n12923), .A2(n1489), .Y(n1481) );
  OR2X1_RVT U1448 ( .A1(n1244), .A2(n1490), .Y(n1480) );
  AND4X1_RVT U1449 ( .A1(n1491), .A2(n1492), .A3(n1493), .A4(n1494), .Y(n1406)
         );
  AND2X1_RVT U1450 ( .A1(n1495), .A2(n1496), .Y(n1494) );
  OR2X1_RVT U1451 ( .A1(n12609), .A2(n1497), .Y(n1496) );
  AND2X1_RVT U1452 ( .A1(n1498), .A2(n1499), .Y(n1495) );
  OR2X1_RVT U1453 ( .A1(n1140), .A2(n1150), .Y(n1499) );
  OR2X1_RVT U1454 ( .A1(n12630), .A2(n1200), .Y(n1150) );
  OR2X1_RVT U1455 ( .A1(n12616), .A2(n1500), .Y(n1498) );
  OR2X1_RVT U1456 ( .A1(n1121), .A2(n1114), .Y(n1493) );
  OR2X1_RVT U1457 ( .A1(n1207), .A2(n1501), .Y(n1114) );
  OR2X1_RVT U1458 ( .A1(n12919), .A2(n1502), .Y(n1492) );
  OR2X1_RVT U1459 ( .A1(n12628), .A2(n1241), .Y(n1491) );
  OR2X1_RVT U1460 ( .A1(n12910), .A2(n1422), .Y(n1241) );
  AND4X1_RVT U1461 ( .A1(n1504), .A2(n1505), .A3(n1506), .A4(n1507), .Y(n1503)
         );
  AND4X1_RVT U1462 ( .A1(n1508), .A2(n1509), .A3(n1510), .A4(n1511), .Y(n1507)
         );
  OR2X1_RVT U1463 ( .A1(n19), .A2(n1512), .Y(n1511) );
  OR2X1_RVT U1464 ( .A1(n1513), .A2(n12641), .Y(n1512) );
  AND2X1_RVT U1465 ( .A1(n12630), .A2(n1160), .Y(n1513) );
  AND2X1_RVT U1466 ( .A1(n1075), .A2(n1514), .Y(n1510) );
  OR2X1_RVT U1467 ( .A1(n12619), .A2(n1515), .Y(n1075) );
  OR2X1_RVT U1468 ( .A1(n19), .A2(n1154), .Y(n1515) );
  OR2X1_RVT U1469 ( .A1(n1516), .A2(n1083), .Y(n1509) );
  AND2X1_RVT U1470 ( .A1(n1517), .A2(n1518), .Y(n1516) );
  AND2X1_RVT U1471 ( .A1(n1519), .A2(n1520), .Y(n1508) );
  OR2X1_RVT U1472 ( .A1(n1521), .A2(n1522), .Y(n1520) );
  AND2X1_RVT U1473 ( .A1(n1523), .A2(n1164), .Y(n1521) );
  OR2X1_RVT U1474 ( .A1(n1524), .A2(n1155), .Y(n1519) );
  AND2X1_RVT U1475 ( .A1(n1459), .A2(n1174), .Y(n1524) );
  OR2X1_RVT U1476 ( .A1(n12617), .A2(n1525), .Y(n1459) );
  OR2X1_RVT U1477 ( .A1(n12925), .A2(n12627), .Y(n1525) );
  AND4X1_RVT U1478 ( .A1(n1526), .A2(n1527), .A3(n1528), .A4(n1529), .Y(n1506)
         );
  OR2X1_RVT U1479 ( .A1(n1530), .A2(n12915), .Y(n1529) );
  AND2X1_RVT U1480 ( .A1(n1223), .A2(n1531), .Y(n1530) );
  OR2X1_RVT U1481 ( .A1(n12923), .A2(n1268), .Y(n1223) );
  AND2X1_RVT U1482 ( .A1(n1532), .A2(n1533), .Y(n1528) );
  OR2X1_RVT U1483 ( .A1(n1534), .A2(n12913), .Y(n1533) );
  AND2X1_RVT U1484 ( .A1(n1535), .A2(n1536), .Y(n1534) );
  OR2X1_RVT U1485 ( .A1(n1118), .A2(n1479), .Y(n1536) );
  OR2X1_RVT U1486 ( .A1(n1537), .A2(n12911), .Y(n1532) );
  AND2X1_RVT U1487 ( .A1(n1538), .A2(n1539), .Y(n1537) );
  OR2X1_RVT U1488 ( .A1(n1540), .A2(n12630), .Y(n1527) );
  AND2X1_RVT U1489 ( .A1(n1541), .A2(n1542), .Y(n1540) );
  AND2X1_RVT U1490 ( .A1(n1543), .A2(n1544), .Y(n1541) );
  AND2X1_RVT U1491 ( .A1(n1545), .A2(n1546), .Y(n1526) );
  OR2X1_RVT U1492 ( .A1(n1547), .A2(n1463), .Y(n1546) );
  AND2X1_RVT U1493 ( .A1(n1548), .A2(n1175), .Y(n1547) );
  AND2X1_RVT U1494 ( .A1(n1549), .A2(n1550), .Y(n1548) );
  OR2X1_RVT U1495 ( .A1(n1551), .A2(n12633), .Y(n1545) );
  AND2X1_RVT U1496 ( .A1(n1552), .A2(n1553), .Y(n1551) );
  OR2X1_RVT U1497 ( .A1(n12922), .A2(n12635), .Y(n1553) );
  AND2X1_RVT U1498 ( .A1(n1164), .A2(n1554), .Y(n1552) );
  AND4X1_RVT U1499 ( .A1(n1555), .A2(n1556), .A3(n1557), .A4(n1558), .Y(n1505)
         );
  AND2X1_RVT U1500 ( .A1(n1559), .A2(n1560), .Y(n1558) );
  OR2X1_RVT U1501 ( .A1(n1157), .A2(n1231), .Y(n1560) );
  OR2X1_RVT U1502 ( .A1(n12917), .A2(n1164), .Y(n1231) );
  AND2X1_RVT U1503 ( .A1(n1561), .A2(n1562), .Y(n1559) );
  OR2X1_RVT U1504 ( .A1(n1428), .A2(n1123), .Y(n1562) );
  OR2X1_RVT U1505 ( .A1(n12924), .A2(n12626), .Y(n1123) );
  OR2X1_RVT U1506 ( .A1(n1207), .A2(n1257), .Y(n1561) );
  OR2X1_RVT U1507 ( .A1(n12912), .A2(n1563), .Y(n1257) );
  OR2X1_RVT U1508 ( .A1(n1564), .A2(n12609), .Y(n1557) );
  AND4X1_RVT U1509 ( .A1(n1565), .A2(n1566), .A3(n1567), .A4(n1568), .Y(n1564)
         );
  OR2X1_RVT U1510 ( .A1(n1501), .A2(n1155), .Y(n1567) );
  OR2X1_RVT U1511 ( .A1(n1569), .A2(n1152), .Y(n1566) );
  OR2X1_RVT U1512 ( .A1(n12921), .A2(n1107), .Y(n1565) );
  OR2X1_RVT U1513 ( .A1(n1570), .A2(n12610), .Y(n1556) );
  AND2X1_RVT U1514 ( .A1(n1571), .A2(n1572), .Y(n1570) );
  OR2X1_RVT U1515 ( .A1(n1501), .A2(n1107), .Y(n1572) );
  AND2X1_RVT U1516 ( .A1(n1573), .A2(n1502), .Y(n1571) );
  OR2X1_RVT U1517 ( .A1(n1155), .A2(n1574), .Y(n1502) );
  OR2X1_RVT U1518 ( .A1(n12912), .A2(n12924), .Y(n1574) );
  OR2X1_RVT U1519 ( .A1(n1575), .A2(n12617), .Y(n1555) );
  AND4X1_RVT U1520 ( .A1(n1576), .A2(n1489), .A3(n1179), .A4(n1151), .Y(n1575)
         );
  OR2X1_RVT U1521 ( .A1(n1176), .A2(n1577), .Y(n1151) );
  OR2X1_RVT U1522 ( .A1(n12914), .A2(n1113), .Y(n1577) );
  OR2X1_RVT U1523 ( .A1(n1238), .A2(n1272), .Y(n1179) );
  OR2X1_RVT U1524 ( .A1(n1157), .A2(n1578), .Y(n1489) );
  OR2X1_RVT U1525 ( .A1(n12641), .A2(n12610), .Y(n1578) );
  OR2X1_RVT U1526 ( .A1(n1116), .A2(n1579), .Y(n1576) );
  OR2X1_RVT U1527 ( .A1(n1580), .A2(n12615), .Y(n1579) );
  AND4X1_RVT U1528 ( .A1(n1581), .A2(n1582), .A3(n1583), .A4(n1584), .Y(n1504)
         );
  AND2X1_RVT U1529 ( .A1(n1585), .A2(n1586), .Y(n1584) );
  AND2X1_RVT U1530 ( .A1(n1587), .A2(n1588), .Y(n1585) );
  OR2X1_RVT U1531 ( .A1(n1148), .A2(n1542), .Y(n1588) );
  OR2X1_RVT U1532 ( .A1(n1160), .A2(n1589), .Y(n1542) );
  OR2X1_RVT U1533 ( .A1(n12913), .A2(n12915), .Y(n1589) );
  OR2X1_RVT U1534 ( .A1(n12920), .A2(n1590), .Y(n1587) );
  OR2X1_RVT U1535 ( .A1(n12626), .A2(n1591), .Y(n1583) );
  OR2X1_RVT U1536 ( .A1(n12923), .A2(n1592), .Y(n1582) );
  OR2X1_RVT U1537 ( .A1(n1160), .A2(n1593), .Y(n1581) );
  AND4X1_RVT U1538 ( .A1(n1595), .A2(n1596), .A3(n1597), .A4(n1598), .Y(n1594)
         );
  AND4X1_RVT U1539 ( .A1(n1599), .A2(n1600), .A3(n1601), .A4(n1602), .Y(n1598)
         );
  AND4X1_RVT U1540 ( .A1(n1603), .A2(n1604), .A3(n1077), .A4(n1605), .Y(n1602)
         );
  OR2X1_RVT U1541 ( .A1(n1218), .A2(n1606), .Y(n1077) );
  OR2X1_RVT U1542 ( .A1(n1428), .A2(n11), .Y(n1606) );
  OR2X1_RVT U1543 ( .A1(n1081), .A2(n1607), .Y(n1604) );
  OR2X1_RVT U1544 ( .A1(n12918), .A2(n12921), .Y(n1607) );
  OR2X1_RVT U1545 ( .A1(n1463), .A2(n1608), .Y(n1603) );
  OR2X1_RVT U1546 ( .A1(n1609), .A2(n1118), .Y(n1608) );
  AND2X1_RVT U1547 ( .A1(n12630), .A2(n1218), .Y(n1609) );
  OR2X1_RVT U1548 ( .A1(n1610), .A2(n12636), .Y(n1601) );
  AND2X1_RVT U1549 ( .A1(n1478), .A2(n1550), .Y(n1610) );
  OR2X1_RVT U1550 ( .A1(n11), .A2(n1611), .Y(n1550) );
  OR2X1_RVT U1551 ( .A1(n12609), .A2(n12917), .Y(n1611) );
  OR2X1_RVT U1552 ( .A1(n1148), .A2(n1612), .Y(n1478) );
  OR2X1_RVT U1553 ( .A1(n12915), .A2(n1140), .Y(n1612) );
  OR2X1_RVT U1554 ( .A1(n1613), .A2(n1098), .Y(n1600) );
  AND2X1_RVT U1555 ( .A1(n1614), .A2(n1422), .Y(n1613) );
  OR2X1_RVT U1556 ( .A1(n1204), .A2(n1198), .Y(n1599) );
  AND4X1_RVT U1557 ( .A1(n1615), .A2(n1616), .A3(n1617), .A4(n1618), .Y(n1597)
         );
  AND2X1_RVT U1558 ( .A1(n1619), .A2(n1620), .Y(n1618) );
  OR2X1_RVT U1559 ( .A1(n1621), .A2(n12630), .Y(n1620) );
  AND2X1_RVT U1560 ( .A1(n1622), .A2(n1171), .Y(n1621) );
  AND2X1_RVT U1561 ( .A1(n1623), .A2(n1624), .Y(n1619) );
  OR2X1_RVT U1562 ( .A1(n1625), .A2(n1154), .Y(n1624) );
  AND2X1_RVT U1563 ( .A1(n1125), .A2(n1097), .Y(n1625) );
  OR2X1_RVT U1564 ( .A1(n12923), .A2(n1196), .Y(n1125) );
  OR2X1_RVT U1565 ( .A1(n1626), .A2(n1207), .Y(n1623) );
  AND2X1_RVT U1566 ( .A1(n1518), .A2(n1627), .Y(n1626) );
  OR2X1_RVT U1567 ( .A1(n12924), .A2(n1235), .Y(n1518) );
  OR2X1_RVT U1568 ( .A1(n1628), .A2(n12915), .Y(n1617) );
  AND2X1_RVT U1569 ( .A1(n1102), .A2(n1629), .Y(n1628) );
  OR2X1_RVT U1570 ( .A1(n1238), .A2(n1162), .Y(n1629) );
  OR2X1_RVT U1571 ( .A1(n1141), .A2(n1463), .Y(n1102) );
  OR2X1_RVT U1572 ( .A1(n1630), .A2(n9), .Y(n1616) );
  AND2X1_RVT U1573 ( .A1(n1152), .A2(n1631), .Y(n1630) );
  OR2X1_RVT U1574 ( .A1(n1632), .A2(n12614), .Y(n1631) );
  AND2X1_RVT U1575 ( .A1(n1633), .A2(n1634), .Y(n1632) );
  OR2X1_RVT U1576 ( .A1(n12916), .A2(n1135), .Y(n1634) );
  OR2X1_RVT U1577 ( .A1(n12641), .A2(n1238), .Y(n1152) );
  OR2X1_RVT U1578 ( .A1(n1635), .A2(n1222), .Y(n1615) );
  AND2X1_RVT U1579 ( .A1(n1155), .A2(n1200), .Y(n1635) );
  OR2X1_RVT U1580 ( .A1(n12912), .A2(n1083), .Y(n1200) );
  AND4X1_RVT U1581 ( .A1(n1636), .A2(n1637), .A3(n1638), .A4(n1639), .Y(n1596)
         );
  AND4X1_RVT U1582 ( .A1(n1640), .A2(n1641), .A3(n1642), .A4(n1643), .Y(n1639)
         );
  OR2X1_RVT U1583 ( .A1(n1644), .A2(n12923), .Y(n1643) );
  AND2X1_RVT U1584 ( .A1(n1258), .A2(n1645), .Y(n1644) );
  OR2X1_RVT U1585 ( .A1(n12638), .A2(n1107), .Y(n1645) );
  OR2X1_RVT U1586 ( .A1(n1646), .A2(n1100), .Y(n1642) );
  AND2X1_RVT U1587 ( .A1(n1647), .A2(n1648), .Y(n1646) );
  OR2X1_RVT U1588 ( .A1(n1649), .A2(n1135), .Y(n1648) );
  AND2X1_RVT U1589 ( .A1(n1160), .A2(n1148), .Y(n1649) );
  AND2X1_RVT U1590 ( .A1(n1162), .A2(n1523), .Y(n1647) );
  OR2X1_RVT U1591 ( .A1(n12639), .A2(n1419), .Y(n1523) );
  OR2X1_RVT U1592 ( .A1(n1650), .A2(n12628), .Y(n1641) );
  AND2X1_RVT U1593 ( .A1(n1651), .A2(n1652), .Y(n1650) );
  OR2X1_RVT U1594 ( .A1(n1148), .A2(n1653), .Y(n1652) );
  AND2X1_RVT U1595 ( .A1(n1230), .A2(n1543), .Y(n1651) );
  OR2X1_RVT U1596 ( .A1(n1140), .A2(n1434), .Y(n1543) );
  OR2X1_RVT U1597 ( .A1(n1113), .A2(n1654), .Y(n1230) );
  OR2X1_RVT U1598 ( .A1(n1655), .A2(n1083), .Y(n1640) );
  AND4X1_RVT U1599 ( .A1(n1656), .A2(n1657), .A3(n1658), .A4(n1591), .Y(n1655)
         );
  OR2X1_RVT U1600 ( .A1(n1176), .A2(n1659), .Y(n1591) );
  OR2X1_RVT U1601 ( .A1(n12609), .A2(n1140), .Y(n1659) );
  OR2X1_RVT U1602 ( .A1(n12920), .A2(n1501), .Y(n1657) );
  OR2X1_RVT U1603 ( .A1(n1141), .A2(n1238), .Y(n1656) );
  OR2X1_RVT U1604 ( .A1(n1428), .A2(n1470), .Y(n1638) );
  OR2X1_RVT U1605 ( .A1(n1660), .A2(n12612), .Y(n1637) );
  AND4X1_RVT U1606 ( .A1(n1661), .A2(n1662), .A3(n1185), .A4(n1283), .Y(n1660)
         );
  OR2X1_RVT U1607 ( .A1(n1107), .A2(n1272), .Y(n1283) );
  OR2X1_RVT U1608 ( .A1(n12920), .A2(n9), .Y(n1272) );
  OR2X1_RVT U1609 ( .A1(n1100), .A2(n1164), .Y(n1185) );
  OR2X1_RVT U1610 ( .A1(n12912), .A2(n1654), .Y(n1636) );
  AND4X1_RVT U1611 ( .A1(n1663), .A2(n1664), .A3(n1665), .A4(n1666), .Y(n1595)
         );
  OR2X1_RVT U1612 ( .A1(n12617), .A2(n1667), .Y(n1666) );
  AND2X1_RVT U1613 ( .A1(n1668), .A2(n1669), .Y(n1665) );
  OR2X1_RVT U1614 ( .A1(n12638), .A2(n1422), .Y(n1669) );
  OR2X1_RVT U1615 ( .A1(n1090), .A2(n1164), .Y(n1668) );
  OR2X1_RVT U1616 ( .A1(n11), .A2(n1121), .Y(n1164) );
  OR2X1_RVT U1617 ( .A1(n12641), .A2(n1282), .Y(n1664) );
  OR2X1_RVT U1618 ( .A1(n1157), .A2(n1670), .Y(n1282) );
  AND2X1_RVT U1619 ( .A1(n1671), .A2(n1672), .Y(n1663) );
  OR2X1_RVT U1620 ( .A1(n12610), .A2(n1673), .Y(n1672) );
  OR2X1_RVT U1621 ( .A1(n1160), .A2(n1109), .Y(n1671) );
  OR2X1_RVT U1622 ( .A1(n1083), .A2(n1487), .Y(n1109) );
  AND4X1_RVT U1623 ( .A1(n1675), .A2(n1676), .A3(n1677), .A4(n1678), .Y(n1674)
         );
  AND4X1_RVT U1624 ( .A1(n1679), .A2(n1680), .A3(n1681), .A4(n1682), .Y(n1678)
         );
  AND4X1_RVT U1625 ( .A1(n1415), .A2(n1605), .A3(n1683), .A4(n1684), .Y(n1682)
         );
  OR2X1_RVT U1626 ( .A1(n1685), .A2(n1686), .Y(n1605) );
  OR2X1_RVT U1627 ( .A1(n1081), .A2(n1470), .Y(n1415) );
  OR2X1_RVT U1628 ( .A1(n12921), .A2(n12626), .Y(n1470) );
  AND4X1_RVT U1629 ( .A1(n1673), .A2(n1539), .A3(n1662), .A4(n1078), .Y(n1681)
         );
  OR2X1_RVT U1630 ( .A1(n1687), .A2(n1268), .Y(n1078) );
  OR2X1_RVT U1631 ( .A1(n1083), .A2(n1688), .Y(n1662) );
  OR2X1_RVT U1632 ( .A1(n1116), .A2(n9), .Y(n1539) );
  OR2X1_RVT U1633 ( .A1(n1107), .A2(n1689), .Y(n1673) );
  OR2X1_RVT U1634 ( .A1(n12616), .A2(n12636), .Y(n1689) );
  AND4X1_RVT U1635 ( .A1(n1690), .A2(n1691), .A3(n1692), .A4(n1693), .Y(n1680)
         );
  OR2X1_RVT U1636 ( .A1(n1479), .A2(n1694), .Y(n1693) );
  OR2X1_RVT U1637 ( .A1(n12636), .A2(n1140), .Y(n1694) );
  OR2X1_RVT U1638 ( .A1(n1269), .A2(n1695), .Y(n1692) );
  OR2X1_RVT U1639 ( .A1(n12922), .A2(n1157), .Y(n1695) );
  OR2X1_RVT U1640 ( .A1(n1614), .A2(n1696), .Y(n1691) );
  OR2X1_RVT U1641 ( .A1(n1697), .A2(n1154), .Y(n1696) );
  OR2X1_RVT U1642 ( .A1(n12633), .A2(n1698), .Y(n1690) );
  OR2X1_RVT U1643 ( .A1(n1699), .A2(n12616), .Y(n1698) );
  AND2X1_RVT U1644 ( .A1(n1487), .A2(n1700), .Y(n1699) );
  AND2X1_RVT U1645 ( .A1(n1701), .A2(n1702), .Y(n1679) );
  OR2X1_RVT U1646 ( .A1(n1703), .A2(n1135), .Y(n1702) );
  AND2X1_RVT U1647 ( .A1(n1704), .A2(n1705), .Y(n1703) );
  OR2X1_RVT U1648 ( .A1(n12615), .A2(n1447), .Y(n1705) );
  OR2X1_RVT U1649 ( .A1(n12619), .A2(n1522), .Y(n1704) );
  AND2X1_RVT U1650 ( .A1(n1706), .A2(n1707), .Y(n1701) );
  OR2X1_RVT U1651 ( .A1(n1708), .A2(n1174), .Y(n1707) );
  AND2X1_RVT U1652 ( .A1(n1709), .A2(n1710), .Y(n1708) );
  OR2X1_RVT U1653 ( .A1(n12622), .A2(n19), .Y(n1710) );
  NAND2X1_RVT U1654 ( .A1(n1157), .A2(n12914), .Y(n1709) );
  OR2X1_RVT U1655 ( .A1(n1711), .A2(n11), .Y(n1706) );
  AND2X1_RVT U1656 ( .A1(n1500), .A2(n1258), .Y(n1711) );
  OR2X1_RVT U1657 ( .A1(n1107), .A2(n1712), .Y(n1258) );
  OR2X1_RVT U1658 ( .A1(n12925), .A2(n12611), .Y(n1712) );
  AND4X1_RVT U1659 ( .A1(n1275), .A2(n1713), .A3(n1586), .A4(n1714), .Y(n1677)
         );
  AND4X1_RVT U1660 ( .A1(n1715), .A2(n1716), .A3(n1717), .A4(n1718), .Y(n1714)
         );
  OR2X1_RVT U1661 ( .A1(n1238), .A2(n1159), .Y(n1718) );
  OR2X1_RVT U1662 ( .A1(n1176), .A2(n1205), .Y(n1717) );
  OR2X1_RVT U1663 ( .A1(n12913), .A2(n1549), .Y(n1716) );
  OR2X1_RVT U1664 ( .A1(n1154), .A2(n1136), .Y(n1549) );
  OR2X1_RVT U1665 ( .A1(n12921), .A2(n1218), .Y(n1136) );
  OR2X1_RVT U1666 ( .A1(n12625), .A2(n1259), .Y(n1715) );
  OR2X1_RVT U1667 ( .A1(n1140), .A2(n1487), .Y(n1259) );
  OR2X1_RVT U1668 ( .A1(n12609), .A2(n1463), .Y(n1487) );
  AND2X1_RVT U1669 ( .A1(n1719), .A2(n1720), .Y(n1586) );
  OR2X1_RVT U1670 ( .A1(n1721), .A2(n1207), .Y(n1720) );
  OR2X1_RVT U1671 ( .A1(n12635), .A2(n11), .Y(n1721) );
  OR2X1_RVT U1672 ( .A1(n1722), .A2(n1090), .Y(n1719) );
  OR2X1_RVT U1673 ( .A1(n12912), .A2(n1207), .Y(n1090) );
  OR2X1_RVT U1674 ( .A1(n1104), .A2(n1154), .Y(n1722) );
  OR2X1_RVT U1675 ( .A1(n12617), .A2(n1592), .Y(n1713) );
  AND2X1_RVT U1676 ( .A1(n1723), .A2(n1724), .Y(n1275) );
  OR2X1_RVT U1677 ( .A1(n1158), .A2(n1196), .Y(n1724) );
  OR2X1_RVT U1678 ( .A1(n1725), .A2(n1726), .Y(n1723) );
  AND4X1_RVT U1679 ( .A1(n1727), .A2(n1728), .A3(n1729), .A4(n1730), .Y(n1676)
         );
  OR2X1_RVT U1680 ( .A1(n1731), .A2(n1463), .Y(n1730) );
  AND2X1_RVT U1681 ( .A1(n1732), .A2(n1472), .Y(n1731) );
  OR2X1_RVT U1682 ( .A1(n12623), .A2(n1688), .Y(n1472) );
  OR2X1_RVT U1683 ( .A1(n1733), .A2(n12918), .Y(n1729) );
  AND2X1_RVT U1684 ( .A1(n1281), .A2(n1246), .Y(n1733) );
  OR2X1_RVT U1685 ( .A1(n12912), .A2(n1222), .Y(n1246) );
  OR2X1_RVT U1686 ( .A1(n1734), .A2(n1420), .Y(n1728) );
  AND2X1_RVT U1687 ( .A1(n1735), .A2(n1736), .Y(n1734) );
  OR2X1_RVT U1688 ( .A1(n12612), .A2(n1160), .Y(n1736) );
  AND2X1_RVT U1689 ( .A1(n1737), .A2(n1198), .Y(n1735) );
  OR2X1_RVT U1690 ( .A1(n9), .A2(n1157), .Y(n1737) );
  OR2X1_RVT U1691 ( .A1(n1738), .A2(n1098), .Y(n1727) );
  AND2X1_RVT U1692 ( .A1(n1739), .A2(n1740), .Y(n1738) );
  NAND2X1_RVT U1693 ( .A1(n1083), .A2(n1580), .Y(n1740) );
  AND2X1_RVT U1694 ( .A1(n1741), .A2(n1430), .Y(n1739) );
  OR2X1_RVT U1695 ( .A1(n1244), .A2(n1688), .Y(n1430) );
  OR2X1_RVT U1696 ( .A1(n12632), .A2(n1742), .Y(n1741) );
  AND4X1_RVT U1697 ( .A1(n1743), .A2(n1744), .A3(n1745), .A4(n1746), .Y(n1675)
         );
  OR2X1_RVT U1698 ( .A1(n1747), .A2(n1121), .Y(n1746) );
  AND2X1_RVT U1699 ( .A1(n1748), .A2(n1262), .Y(n1747) );
  AND2X1_RVT U1700 ( .A1(n1749), .A2(n1284), .Y(n1748) );
  OR2X1_RVT U1701 ( .A1(n11), .A2(n1726), .Y(n1284) );
  OR2X1_RVT U1702 ( .A1(n12611), .A2(n1218), .Y(n1726) );
  OR2X1_RVT U1703 ( .A1(n1750), .A2(n12628), .Y(n1745) );
  AND2X1_RVT U1704 ( .A1(n1751), .A2(n1752), .Y(n1750) );
  OR2X1_RVT U1705 ( .A1(n1753), .A2(n12910), .Y(n1752) );
  AND2X1_RVT U1706 ( .A1(n1754), .A2(n1755), .Y(n1753) );
  OR2X1_RVT U1707 ( .A1(n12610), .A2(n1614), .Y(n1755) );
  OR2X1_RVT U1708 ( .A1(n12917), .A2(n1141), .Y(n1754) );
  AND2X1_RVT U1709 ( .A1(n1756), .A2(n1757), .Y(n1751) );
  OR2X1_RVT U1710 ( .A1(n1107), .A2(n1758), .Y(n1756) );
  OR2X1_RVT U1711 ( .A1(n1759), .A2(n1141), .Y(n1744) );
  AND4X1_RVT U1712 ( .A1(n1760), .A2(n1761), .A3(n1762), .A4(n1107), .Y(n1759)
         );
  OR2X1_RVT U1713 ( .A1(n12918), .A2(n1157), .Y(n1762) );
  OR2X1_RVT U1714 ( .A1(n12622), .A2(n1176), .Y(n1761) );
  OR2X1_RVT U1715 ( .A1(n1229), .A2(n1207), .Y(n1760) );
  OR2X1_RVT U1716 ( .A1(n1763), .A2(n1083), .Y(n1743) );
  AND4X1_RVT U1717 ( .A1(n1627), .A2(n1764), .A3(n1425), .A4(n1222), .Y(n1763)
         );
  OR2X1_RVT U1718 ( .A1(n1176), .A2(n1758), .Y(n1425) );
  OR2X1_RVT U1719 ( .A1(n1463), .A2(n1670), .Y(n1764) );
  OR2X1_RVT U1720 ( .A1(n12616), .A2(n1428), .Y(n1627) );
  AND4X1_RVT U1721 ( .A1(n1766), .A2(n1767), .A3(n1768), .A4(n1769), .Y(n1765)
         );
  AND4X1_RVT U1722 ( .A1(n1159), .A2(n1514), .A3(n1770), .A4(n1771), .Y(n1769)
         );
  AND4X1_RVT U1723 ( .A1(n1593), .A2(n1538), .A3(n1683), .A4(n1684), .Y(n1771)
         );
  OR2X1_RVT U1724 ( .A1(n1686), .A2(n1080), .Y(n1684) );
  OR2X1_RVT U1725 ( .A1(n12916), .A2(n1198), .Y(n1080) );
  OR2X1_RVT U1726 ( .A1(n1097), .A2(n1725), .Y(n1683) );
  OR2X1_RVT U1727 ( .A1(n12921), .A2(n12630), .Y(n1725) );
  OR2X1_RVT U1728 ( .A1(n12910), .A2(n1218), .Y(n1097) );
  OR2X1_RVT U1729 ( .A1(n12922), .A2(n1116), .Y(n1538) );
  OR2X1_RVT U1730 ( .A1(n12639), .A2(n12623), .Y(n1116) );
  OR2X1_RVT U1731 ( .A1(n1238), .A2(n1772), .Y(n1593) );
  OR2X1_RVT U1732 ( .A1(n12630), .A2(n1142), .Y(n1772) );
  OR2X1_RVT U1733 ( .A1(n1140), .A2(n1773), .Y(n1770) );
  OR2X1_RVT U1734 ( .A1(n1268), .A2(n12621), .Y(n1773) );
  OR2X1_RVT U1735 ( .A1(n1207), .A2(n1774), .Y(n1514) );
  OR2X1_RVT U1736 ( .A1(n1141), .A2(n12628), .Y(n1774) );
  OR2X1_RVT U1737 ( .A1(n12914), .A2(n1685), .Y(n1159) );
  OR2X1_RVT U1738 ( .A1(n12623), .A2(n1158), .Y(n1685) );
  AND4X1_RVT U1739 ( .A1(n1775), .A2(n1776), .A3(n1777), .A4(n1778), .Y(n1768)
         );
  AND4X1_RVT U1740 ( .A1(n1779), .A2(n1780), .A3(n1781), .A4(n1782), .Y(n1778)
         );
  OR2X1_RVT U1741 ( .A1(n1174), .A2(n1783), .Y(n1782) );
  OR2X1_RVT U1742 ( .A1(n12612), .A2(n1244), .Y(n1783) );
  OR2X1_RVT U1743 ( .A1(n1157), .A2(n1784), .Y(n1781) );
  OR2X1_RVT U1744 ( .A1(n1785), .A2(n1121), .Y(n1784) );
  AND2X1_RVT U1745 ( .A1(n1100), .A2(n1160), .Y(n1785) );
  OR2X1_RVT U1746 ( .A1(n1786), .A2(n1787), .Y(n1780) );
  AND2X1_RVT U1747 ( .A1(n1434), .A2(n1271), .Y(n1786) );
  OR2X1_RVT U1748 ( .A1(n12915), .A2(n19), .Y(n1271) );
  OR2X1_RVT U1749 ( .A1(n12911), .A2(n12633), .Y(n1434) );
  OR2X1_RVT U1750 ( .A1(n1788), .A2(n1155), .Y(n1779) );
  AND2X1_RVT U1751 ( .A1(n1670), .A2(n1789), .Y(n1788) );
  OR2X1_RVT U1752 ( .A1(n12913), .A2(n11), .Y(n1789) );
  OR2X1_RVT U1753 ( .A1(n1790), .A2(n12635), .Y(n1777) );
  AND2X1_RVT U1754 ( .A1(n1661), .A2(n1791), .Y(n1790) );
  OR2X1_RVT U1755 ( .A1(n1148), .A2(n1614), .Y(n1791) );
  OR2X1_RVT U1756 ( .A1(n12616), .A2(n1479), .Y(n1661) );
  OR2X1_RVT U1757 ( .A1(n12917), .A2(n1148), .Y(n1479) );
  OR2X1_RVT U1758 ( .A1(n1792), .A2(n1428), .Y(n1776) );
  AND2X1_RVT U1759 ( .A1(n1262), .A2(n1653), .Y(n1792) );
  OR2X1_RVT U1760 ( .A1(n1118), .A2(n1207), .Y(n1262) );
  OR2X1_RVT U1761 ( .A1(n1793), .A2(n1198), .Y(n1775) );
  AND2X1_RVT U1762 ( .A1(n1161), .A2(n1163), .Y(n1793) );
  AND4X1_RVT U1763 ( .A1(n1794), .A2(n1795), .A3(n1796), .A4(n1797), .Y(n1767)
         );
  AND4X1_RVT U1764 ( .A1(n1798), .A2(n1799), .A3(n1800), .A4(n1801), .Y(n1797)
         );
  OR2X1_RVT U1765 ( .A1(n1802), .A2(n12619), .Y(n1801) );
  AND2X1_RVT U1766 ( .A1(n1089), .A2(n1500), .Y(n1802) );
  OR2X1_RVT U1767 ( .A1(n1238), .A2(n1269), .Y(n1500) );
  OR2X1_RVT U1768 ( .A1(n12622), .A2(n1121), .Y(n1269) );
  OR2X1_RVT U1769 ( .A1(n12626), .A2(n1803), .Y(n1089) );
  OR2X1_RVT U1770 ( .A1(n12609), .A2(n12615), .Y(n1803) );
  OR2X1_RVT U1771 ( .A1(n1804), .A2(n12633), .Y(n1800) );
  AND2X1_RVT U1772 ( .A1(n1517), .A2(n1805), .Y(n1804) );
  OR2X1_RVT U1773 ( .A1(n12638), .A2(n9), .Y(n1805) );
  OR2X1_RVT U1774 ( .A1(n12636), .A2(n1205), .Y(n1517) );
  OR2X1_RVT U1775 ( .A1(n1806), .A2(n12614), .Y(n1799) );
  AND2X1_RVT U1776 ( .A1(n1535), .A2(n1807), .Y(n1806) );
  OR2X1_RVT U1777 ( .A1(n12639), .A2(n1141), .Y(n1807) );
  OR2X1_RVT U1778 ( .A1(n1083), .A2(n1808), .Y(n1535) );
  OR2X1_RVT U1779 ( .A1(n1809), .A2(n1142), .Y(n1798) );
  AND2X1_RVT U1780 ( .A1(n1810), .A2(n1811), .Y(n1809) );
  OR2X1_RVT U1781 ( .A1(n1198), .A2(n12636), .Y(n1811) );
  AND2X1_RVT U1782 ( .A1(n1812), .A2(n1174), .Y(n1810) );
  OR2X1_RVT U1783 ( .A1(n1160), .A2(n1121), .Y(n1174) );
  OR2X1_RVT U1784 ( .A1(n12611), .A2(n1205), .Y(n1812) );
  OR2X1_RVT U1785 ( .A1(n12925), .A2(n1160), .Y(n1205) );
  OR2X1_RVT U1786 ( .A1(n1813), .A2(n1218), .Y(n1796) );
  AND4X1_RVT U1787 ( .A1(n1814), .A2(n1815), .A3(n1490), .A4(n1281), .Y(n1813)
         );
  OR2X1_RVT U1788 ( .A1(n1463), .A2(n1563), .Y(n1281) );
  OR2X1_RVT U1789 ( .A1(n1176), .A2(n1742), .Y(n1490) );
  OR2X1_RVT U1790 ( .A1(n12617), .A2(n12610), .Y(n1742) );
  OR2X1_RVT U1791 ( .A1(n11), .A2(n1098), .Y(n1815) );
  OR2X1_RVT U1792 ( .A1(n9), .A2(n12636), .Y(n1814) );
  OR2X1_RVT U1793 ( .A1(n1816), .A2(n1154), .Y(n1795) );
  AND2X1_RVT U1794 ( .A1(n1817), .A2(n1175), .Y(n1816) );
  AND2X1_RVT U1795 ( .A1(n1749), .A2(n1544), .Y(n1817) );
  OR2X1_RVT U1796 ( .A1(n1818), .A2(n12922), .Y(n1544) );
  AND2X1_RVT U1797 ( .A1(n1196), .A2(n1819), .Y(n1818) );
  OR2X1_RVT U1798 ( .A1(n12614), .A2(n1083), .Y(n1819) );
  OR2X1_RVT U1799 ( .A1(n1244), .A2(n1501), .Y(n1749) );
  OR2X1_RVT U1800 ( .A1(n1229), .A2(n1118), .Y(n1501) );
  OR2X1_RVT U1801 ( .A1(n1820), .A2(n1222), .Y(n1794) );
  AND2X1_RVT U1802 ( .A1(n1821), .A2(n12622), .Y(n1820) );
  AND2X1_RVT U1803 ( .A1(n1822), .A2(n1522), .Y(n1821) );
  OR2X1_RVT U1804 ( .A1(n1244), .A2(n1463), .Y(n1822) );
  AND4X1_RVT U1805 ( .A1(n1823), .A2(n1824), .A3(n1825), .A4(n1826), .Y(n1766)
         );
  AND2X1_RVT U1806 ( .A1(n1827), .A2(n1828), .Y(n1826) );
  OR2X1_RVT U1807 ( .A1(n12918), .A2(n1443), .Y(n1828) );
  OR2X1_RVT U1808 ( .A1(n12630), .A2(n1829), .Y(n1443) );
  OR2X1_RVT U1809 ( .A1(n1140), .A2(n1229), .Y(n1829) );
  AND2X1_RVT U1810 ( .A1(n1830), .A2(n1831), .Y(n1827) );
  OR2X1_RVT U1811 ( .A1(n1113), .A2(n1124), .Y(n1831) );
  OR2X1_RVT U1812 ( .A1(n1157), .A2(n1471), .Y(n1124) );
  OR2X1_RVT U1813 ( .A1(n12914), .A2(n1118), .Y(n1471) );
  OR2X1_RVT U1814 ( .A1(n1160), .A2(n1237), .Y(n1830) );
  OR2X1_RVT U1815 ( .A1(n1148), .A2(n1832), .Y(n1237) );
  OR2X1_RVT U1816 ( .A1(n1148), .A2(n1447), .Y(n1825) );
  OR2X1_RVT U1817 ( .A1(n11), .A2(n12632), .Y(n1447) );
  OR2X1_RVT U1818 ( .A1(n1833), .A2(n1104), .Y(n1824) );
  AND4X1_RVT U1819 ( .A1(n1834), .A2(n1835), .A3(n1836), .A4(n1837), .Y(n1833)
         );
  OR2X1_RVT U1820 ( .A1(n12912), .A2(n1838), .Y(n1836) );
  OR2X1_RVT U1821 ( .A1(n1839), .A2(n12919), .Y(n1838) );
  AND2X1_RVT U1822 ( .A1(n1155), .A2(n1840), .Y(n1839) );
  OR2X1_RVT U1823 ( .A1(n12625), .A2(n1841), .Y(n1835) );
  OR2X1_RVT U1824 ( .A1(n1580), .A2(n1098), .Y(n1841) );
  OR2X1_RVT U1825 ( .A1(n1081), .A2(n1107), .Y(n1834) );
  OR2X1_RVT U1826 ( .A1(n12916), .A2(n1207), .Y(n1107) );
  OR2X1_RVT U1827 ( .A1(n1700), .A2(n1614), .Y(n1823) );
  OR2X1_RVT U1828 ( .A1(n12641), .A2(n1118), .Y(n1614) );
  AND4X1_RVT U1829 ( .A1(n1843), .A2(n1844), .A3(n1845), .A4(n1846), .Y(n1842)
         );
  AND4X1_RVT U1830 ( .A1(n1847), .A2(n1848), .A3(n1849), .A4(n1850), .Y(n1846)
         );
  AND4X1_RVT U1831 ( .A1(n1851), .A2(n1852), .A3(n1853), .A4(n1854), .Y(n1850)
         );
  OR2X1_RVT U1832 ( .A1(n1688), .A2(n1832), .Y(n1854) );
  OR2X1_RVT U1833 ( .A1(n12915), .A2(n12635), .Y(n1832) );
  OR2X1_RVT U1834 ( .A1(n12609), .A2(n12619), .Y(n1688) );
  OR2X1_RVT U1835 ( .A1(n1855), .A2(n1155), .Y(n1853) );
  AND2X1_RVT U1836 ( .A1(n1101), .A2(n1787), .Y(n1855) );
  OR2X1_RVT U1837 ( .A1(n11), .A2(n1856), .Y(n1101) );
  OR2X1_RVT U1838 ( .A1(n12609), .A2(n12912), .Y(n1856) );
  OR2X1_RVT U1839 ( .A1(n1857), .A2(n1083), .Y(n1852) );
  OR2X1_RVT U1840 ( .A1(n12623), .A2(n1244), .Y(n1083) );
  AND2X1_RVT U1841 ( .A1(n1219), .A2(n1858), .Y(n1857) );
  OR2X1_RVT U1842 ( .A1(n1098), .A2(n1419), .Y(n1858) );
  OR2X1_RVT U1843 ( .A1(n12627), .A2(n12615), .Y(n1098) );
  OR2X1_RVT U1844 ( .A1(n1463), .A2(n1859), .Y(n1219) );
  OR2X1_RVT U1845 ( .A1(n12923), .A2(n12630), .Y(n1859) );
  OR2X1_RVT U1846 ( .A1(n1860), .A2(n1142), .Y(n1851) );
  AND2X1_RVT U1847 ( .A1(n1658), .A2(n1861), .Y(n1860) );
  OR2X1_RVT U1848 ( .A1(n1862), .A2(n12912), .Y(n1861) );
  AND2X1_RVT U1849 ( .A1(n1198), .A2(n1670), .Y(n1862) );
  OR2X1_RVT U1850 ( .A1(n12920), .A2(n1160), .Y(n1670) );
  OR2X1_RVT U1851 ( .A1(n12636), .A2(n1863), .Y(n1658) );
  OR2X1_RVT U1852 ( .A1(n12925), .A2(n12921), .Y(n1863) );
  OR2X1_RVT U1853 ( .A1(n1864), .A2(n12614), .Y(n1849) );
  AND2X1_RVT U1854 ( .A1(n1865), .A2(n1866), .Y(n1864) );
  OR2X1_RVT U1855 ( .A1(n1867), .A2(n1244), .Y(n1866) );
  AND2X1_RVT U1856 ( .A1(n1428), .A2(n1868), .Y(n1867) );
  OR2X1_RVT U1857 ( .A1(n1100), .A2(n1222), .Y(n1865) );
  OR2X1_RVT U1858 ( .A1(n12628), .A2(n1158), .Y(n1222) );
  OR2X1_RVT U1859 ( .A1(n1869), .A2(n12921), .Y(n1848) );
  AND2X1_RVT U1860 ( .A1(n1433), .A2(n1592), .Y(n1869) );
  OR2X1_RVT U1861 ( .A1(n12626), .A2(n1870), .Y(n1592) );
  OR2X1_RVT U1862 ( .A1(n1154), .A2(n12615), .Y(n1870) );
  OR2X1_RVT U1863 ( .A1(n1100), .A2(n1700), .Y(n1433) );
  OR2X1_RVT U1864 ( .A1(n12615), .A2(n12630), .Y(n1700) );
  OR2X1_RVT U1865 ( .A1(n1871), .A2(n12612), .Y(n1847) );
  AND2X1_RVT U1866 ( .A1(n1473), .A2(n1872), .Y(n1871) );
  OR2X1_RVT U1867 ( .A1(n1687), .A2(n1148), .Y(n1872) );
  OR2X1_RVT U1868 ( .A1(n1207), .A2(n1808), .Y(n1473) );
  OR2X1_RVT U1869 ( .A1(n12920), .A2(n11), .Y(n1808) );
  AND2X1_RVT U1870 ( .A1(n12616), .A2(n12923), .Y(n1569) );
  AND4X1_RVT U1871 ( .A1(n1873), .A2(n1874), .A3(n1875), .A4(n1876), .Y(n1845)
         );
  AND4X1_RVT U1872 ( .A1(n1877), .A2(n1878), .A3(n1879), .A4(n1880), .Y(n1876)
         );
  OR2X1_RVT U1873 ( .A1(n1881), .A2(n12621), .Y(n1880) );
  AND2X1_RVT U1874 ( .A1(n1460), .A2(n1531), .Y(n1881) );
  OR2X1_RVT U1875 ( .A1(n1157), .A2(n1787), .Y(n1531) );
  OR2X1_RVT U1876 ( .A1(n12923), .A2(n1154), .Y(n1787) );
  OR2X1_RVT U1877 ( .A1(n12910), .A2(n12611), .Y(n1157) );
  OR2X1_RVT U1878 ( .A1(n12612), .A2(n1563), .Y(n1460) );
  OR2X1_RVT U1879 ( .A1(n12616), .A2(n12630), .Y(n1563) );
  OR2X1_RVT U1880 ( .A1(n1882), .A2(n12919), .Y(n1879) );
  AND2X1_RVT U1881 ( .A1(n1622), .A2(n1883), .Y(n1882) );
  OR2X1_RVT U1882 ( .A1(n1580), .A2(n1171), .Y(n1883) );
  OR2X1_RVT U1883 ( .A1(n1463), .A2(n1884), .Y(n1171) );
  OR2X1_RVT U1884 ( .A1(n12641), .A2(n12617), .Y(n1884) );
  OR2X1_RVT U1885 ( .A1(n12625), .A2(n1885), .Y(n1622) );
  OR2X1_RVT U1886 ( .A1(n1463), .A2(n1140), .Y(n1885) );
  OR2X1_RVT U1887 ( .A1(n1886), .A2(n12925), .Y(n1878) );
  AND2X1_RVT U1888 ( .A1(n1568), .A2(n1497), .Y(n1886) );
  OR2X1_RVT U1889 ( .A1(n1160), .A2(n1196), .Y(n1497) );
  OR2X1_RVT U1890 ( .A1(n12917), .A2(n1463), .Y(n1196) );
  OR2X1_RVT U1891 ( .A1(n1687), .A2(n1176), .Y(n1568) );
  OR2X1_RVT U1892 ( .A1(n12622), .A2(n12922), .Y(n1687) );
  OR2X1_RVT U1893 ( .A1(n1887), .A2(n1218), .Y(n1877) );
  AND2X1_RVT U1894 ( .A1(n1888), .A2(n1889), .Y(n1887) );
  OR2X1_RVT U1895 ( .A1(n1140), .A2(n1686), .Y(n1889) );
  OR2X1_RVT U1896 ( .A1(n12919), .A2(n19), .Y(n1686) );
  AND2X1_RVT U1897 ( .A1(n1890), .A2(n1554), .Y(n1888) );
  OR2X1_RVT U1898 ( .A1(n1148), .A2(n1891), .Y(n1554) );
  OR2X1_RVT U1899 ( .A1(n12638), .A2(n12617), .Y(n1891) );
  OR2X1_RVT U1900 ( .A1(n1204), .A2(n1141), .Y(n1875) );
  OR2X1_RVT U1901 ( .A1(n12912), .A2(n1100), .Y(n1204) );
  OR2X1_RVT U1902 ( .A1(n1892), .A2(n1104), .Y(n1874) );
  AND2X1_RVT U1903 ( .A1(n1893), .A2(n1285), .Y(n1892) );
  AND2X1_RVT U1904 ( .A1(n1894), .A2(n1895), .Y(n1285) );
  OR2X1_RVT U1905 ( .A1(n12626), .A2(n1428), .Y(n1895) );
  OR2X1_RVT U1906 ( .A1(n1207), .A2(n1081), .Y(n1894) );
  OR2X1_RVT U1907 ( .A1(n12611), .A2(n1154), .Y(n1081) );
  AND2X1_RVT U1908 ( .A1(n1896), .A2(n1590), .Y(n1893) );
  OR2X1_RVT U1909 ( .A1(n1238), .A2(n1840), .Y(n1590) );
  OR2X1_RVT U1910 ( .A1(n12914), .A2(n9), .Y(n1840) );
  OR2X1_RVT U1911 ( .A1(n1100), .A2(n1267), .Y(n1896) );
  OR2X1_RVT U1912 ( .A1(n12610), .A2(n1897), .Y(n1267) );
  OR2X1_RVT U1913 ( .A1(n12910), .A2(n12639), .Y(n1897) );
  OR2X1_RVT U1914 ( .A1(n1898), .A2(n12910), .Y(n1873) );
  AND4X1_RVT U1915 ( .A1(n1899), .A2(n1900), .A3(n1901), .A4(n1732), .Y(n1898)
         );
  OR2X1_RVT U1916 ( .A1(n1154), .A2(n1653), .Y(n1732) );
  OR2X1_RVT U1917 ( .A1(n12915), .A2(n12921), .Y(n1653) );
  OR2X1_RVT U1918 ( .A1(n1154), .A2(n1902), .Y(n1901) );
  OR2X1_RVT U1919 ( .A1(n12616), .A2(n12621), .Y(n1902) );
  OR2X1_RVT U1920 ( .A1(n12920), .A2(n1113), .Y(n1154) );
  OR2X1_RVT U1921 ( .A1(n1903), .A2(n1235), .Y(n1900) );
  OR2X1_RVT U1922 ( .A1(n12610), .A2(n1079), .Y(n1235) );
  AND2X1_RVT U1923 ( .A1(n1218), .A2(n1904), .Y(n1903) );
  OR2X1_RVT U1924 ( .A1(n12918), .A2(n1118), .Y(n1904) );
  OR2X1_RVT U1925 ( .A1(n12914), .A2(n12621), .Y(n1218) );
  OR2X1_RVT U1926 ( .A1(n12916), .A2(n1868), .Y(n1899) );
  OR2X1_RVT U1927 ( .A1(n12920), .A2(n1158), .Y(n1868) );
  OR2X1_RVT U1928 ( .A1(n1104), .A2(n9), .Y(n1158) );
  AND4X1_RVT U1929 ( .A1(n1905), .A2(n1906), .A3(n1907), .A4(n1908), .Y(n1844)
         );
  AND4X1_RVT U1930 ( .A1(n1909), .A2(n1910), .A3(n1911), .A4(n1912), .Y(n1908)
         );
  OR2X1_RVT U1931 ( .A1(n1176), .A2(n1422), .Y(n1912) );
  OR2X1_RVT U1932 ( .A1(n12623), .A2(n1198), .Y(n1422) );
  OR2X1_RVT U1933 ( .A1(n12627), .A2(n1463), .Y(n1176) );
  OR2X1_RVT U1934 ( .A1(n1163), .A2(n1758), .Y(n1911) );
  OR2X1_RVT U1935 ( .A1(n12924), .A2(n12610), .Y(n1758) );
  OR2X1_RVT U1936 ( .A1(n1229), .A2(n1155), .Y(n1163) );
  OR2X1_RVT U1937 ( .A1(n1148), .A2(n1175), .Y(n1910) );
  OR2X1_RVT U1938 ( .A1(n12619), .A2(n12632), .Y(n1175) );
  OR2X1_RVT U1939 ( .A1(n12609), .A2(n12911), .Y(n1148) );
  OR2X1_RVT U1940 ( .A1(n19), .A2(n1633), .Y(n1909) );
  OR2X1_RVT U1941 ( .A1(n12617), .A2(n1420), .Y(n1633) );
  OR2X1_RVT U1942 ( .A1(n1118), .A2(n1667), .Y(n1907) );
  OR2X1_RVT U1943 ( .A1(n19), .A2(n1913), .Y(n1667) );
  OR2X1_RVT U1944 ( .A1(n12917), .A2(n12630), .Y(n1913) );
  AND2X1_RVT U1945 ( .A1(n12611), .A2(n12614), .Y(n1697) );
  OR2X1_RVT U1946 ( .A1(n1160), .A2(n1108), .Y(n1906) );
  OR2X1_RVT U1947 ( .A1(n12639), .A2(n1914), .Y(n1108) );
  OR2X1_RVT U1948 ( .A1(n12918), .A2(n12910), .Y(n1914) );
  OR2X1_RVT U1949 ( .A1(n12616), .A2(n1140), .Y(n1160) );
  OR2X1_RVT U1950 ( .A1(n1207), .A2(n1890), .Y(n1905) );
  OR2X1_RVT U1951 ( .A1(n12612), .A2(n1162), .Y(n1890) );
  OR2X1_RVT U1952 ( .A1(n12920), .A2(n12921), .Y(n1162) );
  AND4X1_RVT U1953 ( .A1(n1915), .A2(n1273), .A3(n1916), .A4(n1917), .Y(n1843)
         );
  OR2X1_RVT U1954 ( .A1(n12616), .A2(n1837), .Y(n1917) );
  OR2X1_RVT U1955 ( .A1(n12916), .A2(n1268), .Y(n1837) );
  OR2X1_RVT U1956 ( .A1(n12614), .A2(n1428), .Y(n1268) );
  OR2X1_RVT U1957 ( .A1(n12609), .A2(n1135), .Y(n1428) );
  AND2X1_RVT U1958 ( .A1(n1918), .A2(n1919), .Y(n1916) );
  OR2X1_RVT U1959 ( .A1(n12638), .A2(n1757), .Y(n1919) );
  OR2X1_RVT U1960 ( .A1(n1207), .A2(n1419), .Y(n1757) );
  OR2X1_RVT U1961 ( .A1(n12616), .A2(n12610), .Y(n1419) );
  OR2X1_RVT U1962 ( .A1(n12611), .A2(n1096), .Y(n1135) );
  OR2X1_RVT U1963 ( .A1(n12923), .A2(n1488), .Y(n1918) );
  OR2X1_RVT U1964 ( .A1(n12635), .A2(n1522), .Y(n1488) );
  OR2X1_RVT U1965 ( .A1(n12915), .A2(n12910), .Y(n1522) );
  OR2X1_RVT U1966 ( .A1(n12913), .A2(n12627), .Y(n1079) );
  AND2X1_RVT U1967 ( .A1(n1920), .A2(n1921), .Y(n1273) );
  OR2X1_RVT U1968 ( .A1(n1155), .A2(n1141), .Y(n1921) );
  OR2X1_RVT U1969 ( .A1(n12922), .A2(n1113), .Y(n1141) );
  AND2X1_RVT U1970 ( .A1(n1140), .A2(n1104), .Y(n1193) );
  OR2X1_RVT U1971 ( .A1(n12622), .A2(n1207), .Y(n1155) );
  OR2X1_RVT U1972 ( .A1(n12911), .A2(n1244), .Y(n1207) );
  OR2X1_RVT U1973 ( .A1(n1922), .A2(n1198), .Y(n1920) );
  OR2X1_RVT U1974 ( .A1(n12616), .A2(n9), .Y(n1198) );
  AND2X1_RVT U1975 ( .A1(n12924), .A2(n12609), .Y(n1580) );
  OR2X1_RVT U1976 ( .A1(n12615), .A2(n1420), .Y(n1922) );
  OR2X1_RVT U1977 ( .A1(n12920), .A2(n12632), .Y(n1420) );
  AND2X1_RVT U1978 ( .A1(n1923), .A2(n1924), .Y(n1915) );
  OR2X1_RVT U1979 ( .A1(n1121), .A2(n1573), .Y(n1924) );
  OR2X1_RVT U1980 ( .A1(n12617), .A2(n1161), .Y(n1573) );
  OR2X1_RVT U1981 ( .A1(n12632), .A2(n1238), .Y(n1161) );
  OR2X1_RVT U1982 ( .A1(n12612), .A2(n12615), .Y(n1238) );
  OR2X1_RVT U1983 ( .A1(n12917), .A2(n12915), .Y(n1100) );
  OR2X1_RVT U1984 ( .A1(n12925), .A2(n12919), .Y(n1121) );
  XOR2X1_RVT U1985 ( .A1(key[124]), .A2(state[124]), .Y(n1096) );
  OR2X1_RVT U1986 ( .A1(n1113), .A2(n1242), .Y(n1923) );
  OR2X1_RVT U1987 ( .A1(n1463), .A2(n1654), .Y(n1242) );
  OR2X1_RVT U1988 ( .A1(n12619), .A2(n1142), .Y(n1654) );
  OR2X1_RVT U1989 ( .A1(n12918), .A2(n1244), .Y(n1142) );
  XOR2X1_RVT U1990 ( .A1(key[122]), .A2(state[122]), .Y(n1244) );
  XOR2X1_RVT U1991 ( .A1(key[123]), .A2(state[123]), .Y(n1178) );
  OR2X1_RVT U1992 ( .A1(n12923), .A2(n12617), .Y(n1118) );
  XOR2X1_RVT U1993 ( .A1(key[125]), .A2(state[125]), .Y(n1104) );
  XOR2X1_RVT U1994 ( .A1(key[126]), .A2(state[126]), .Y(n1140) );
  OR2X1_RVT U1995 ( .A1(n12913), .A2(n12615), .Y(n1463) );
  XOR2X1_RVT U1996 ( .A1(key[120]), .A2(state[120]), .Y(n1119) );
  XOR2X1_RVT U1997 ( .A1(key[121]), .A2(state[121]), .Y(n1229) );
  XOR2X1_RVT U1998 ( .A1(key[127]), .A2(state[127]), .Y(n1113) );
  AND4X1_RVT U1999 ( .A1(n1926), .A2(n1927), .A3(n1928), .A4(n1929), .Y(n1925)
         );
  AND4X1_RVT U2000 ( .A1(n1930), .A2(n1931), .A3(n1932), .A4(n1933), .Y(n1929)
         );
  AND4X1_RVT U2001 ( .A1(n1934), .A2(n1935), .A3(n1936), .A4(n1937), .Y(n1933)
         );
  OR2X1_RVT U2002 ( .A1(n12603), .A2(n1939), .Y(n1932) );
  OR2X1_RVT U2003 ( .A1(n1940), .A2(n1941), .Y(n1930) );
  OR2X1_RVT U2004 ( .A1(n12907), .A2(n1942), .Y(n1941) );
  AND4X1_RVT U2005 ( .A1(n1943), .A2(n1944), .A3(n1945), .A4(n1946), .Y(n1928)
         );
  OR2X1_RVT U2006 ( .A1(n1947), .A2(n12905), .Y(n1946) );
  AND2X1_RVT U2007 ( .A1(n1948), .A2(n1949), .Y(n1947) );
  AND2X1_RVT U2008 ( .A1(n1950), .A2(n1951), .Y(n1945) );
  OR2X1_RVT U2009 ( .A1(n1952), .A2(n31), .Y(n1951) );
  AND2X1_RVT U2010 ( .A1(n1953), .A2(n1954), .Y(n1952) );
  OR2X1_RVT U2011 ( .A1(n12594), .A2(n1956), .Y(n1954) );
  OR2X1_RVT U2012 ( .A1(n1942), .A2(n1957), .Y(n1953) );
  OR2X1_RVT U2013 ( .A1(n1958), .A2(n12600), .Y(n1950) );
  AND2X1_RVT U2014 ( .A1(n1960), .A2(n1961), .Y(n1958) );
  OR2X1_RVT U2015 ( .A1(n1962), .A2(n1963), .Y(n1944) );
  AND2X1_RVT U2016 ( .A1(n1964), .A2(n1965), .Y(n1962) );
  OR2X1_RVT U2017 ( .A1(n12595), .A2(n1966), .Y(n1965) );
  AND2X1_RVT U2018 ( .A1(n1967), .A2(n1968), .Y(n1964) );
  AND2X1_RVT U2019 ( .A1(n1969), .A2(n1970), .Y(n1943) );
  OR2X1_RVT U2020 ( .A1(n1971), .A2(n12577), .Y(n1970) );
  AND2X1_RVT U2021 ( .A1(n1973), .A2(n1974), .Y(n1971) );
  OR2X1_RVT U2022 ( .A1(n1975), .A2(n1976), .Y(n1974) );
  OR2X1_RVT U2023 ( .A1(n12586), .A2(n12581), .Y(n1976) );
  OR2X1_RVT U2024 ( .A1(n1979), .A2(n1980), .Y(n1969) );
  AND2X1_RVT U2025 ( .A1(n1981), .A2(n1982), .Y(n1979) );
  AND2X1_RVT U2026 ( .A1(n1983), .A2(n1984), .Y(n1981) );
  AND4X1_RVT U2027 ( .A1(n1985), .A2(n1986), .A3(n1987), .A4(n1988), .Y(n1927)
         );
  AND4X1_RVT U2028 ( .A1(n1989), .A2(n1990), .A3(n1991), .A4(n1992), .Y(n1988)
         );
  OR2X1_RVT U2029 ( .A1(n1993), .A2(n12606), .Y(n1992) );
  AND4X1_RVT U2030 ( .A1(n1995), .A2(n1996), .A3(n1997), .A4(n1998), .Y(n1993)
         );
  OR2X1_RVT U2031 ( .A1(n1999), .A2(n1966), .Y(n1998) );
  OR2X1_RVT U2032 ( .A1(n2000), .A2(n12592), .Y(n1997) );
  OR2X1_RVT U2033 ( .A1(n2002), .A2(n12583), .Y(n1991) );
  AND4X1_RVT U2034 ( .A1(n2003), .A2(n2004), .A3(n2005), .A4(n2006), .Y(n2002)
         );
  OR2X1_RVT U2035 ( .A1(n2007), .A2(n2008), .Y(n2006) );
  OR2X1_RVT U2036 ( .A1(n12600), .A2(n12595), .Y(n2008) );
  AND2X1_RVT U2037 ( .A1(n2009), .A2(n2010), .Y(n2005) );
  OR2X1_RVT U2038 ( .A1(n12909), .A2(n2011), .Y(n2004) );
  OR2X1_RVT U2039 ( .A1(n2012), .A2(n2013), .Y(n2003) );
  AND2X1_RVT U2040 ( .A1(n2014), .A2(n2015), .Y(n2012) );
  OR2X1_RVT U2041 ( .A1(n12600), .A2(n2016), .Y(n2015) );
  OR2X1_RVT U2042 ( .A1(n1949), .A2(n2017), .Y(n1990) );
  OR2X1_RVT U2043 ( .A1(n2016), .A2(n2018), .Y(n1989) );
  OR2X1_RVT U2044 ( .A1(n2019), .A2(n2020), .Y(n1987) );
  OR2X1_RVT U2045 ( .A1(n2021), .A2(n2014), .Y(n1986) );
  OR2X1_RVT U2046 ( .A1(n2022), .A2(n2023), .Y(n1985) );
  AND4X1_RVT U2047 ( .A1(n2024), .A2(n2025), .A3(n2026), .A4(n2027), .Y(n1926)
         );
  AND2X1_RVT U2048 ( .A1(n2028), .A2(n2029), .Y(n2027) );
  OR2X1_RVT U2049 ( .A1(n2013), .A2(n2030), .Y(n2029) );
  AND2X1_RVT U2050 ( .A1(n2031), .A2(n2032), .Y(n2028) );
  OR2X1_RVT U2051 ( .A1(n2033), .A2(n1956), .Y(n2032) );
  OR2X1_RVT U2052 ( .A1(n1957), .A2(n2034), .Y(n2031) );
  OR2X1_RVT U2053 ( .A1(n29), .A2(n2035), .Y(n2026) );
  OR2X1_RVT U2054 ( .A1(n2036), .A2(n12590), .Y(n2025) );
  OR2X1_RVT U2055 ( .A1(n12593), .A2(n2038), .Y(n2024) );
  AND4X1_RVT U2056 ( .A1(n2040), .A2(n2041), .A3(n2042), .A4(n2043), .Y(n2039)
         );
  AND4X1_RVT U2057 ( .A1(n2044), .A2(n1935), .A3(n2045), .A4(n2046), .Y(n2043)
         );
  AND4X1_RVT U2058 ( .A1(n2047), .A2(n2048), .A3(n2049), .A4(n2050), .Y(n2046)
         );
  OR2X1_RVT U2059 ( .A1(n1956), .A2(n2051), .Y(n2050) );
  OR2X1_RVT U2060 ( .A1(n2052), .A2(n12605), .Y(n2051) );
  OR2X1_RVT U2061 ( .A1(n1957), .A2(n2053), .Y(n2049) );
  OR2X1_RVT U2062 ( .A1(n29), .A2(n12589), .Y(n2053) );
  OR2X1_RVT U2063 ( .A1(n2054), .A2(n2000), .Y(n2048) );
  AND2X1_RVT U2064 ( .A1(n2011), .A2(n2055), .Y(n2054) );
  OR2X1_RVT U2065 ( .A1(n2056), .A2(n2057), .Y(n2047) );
  AND2X1_RVT U2066 ( .A1(n2058), .A2(n2059), .Y(n2056) );
  AND2X1_RVT U2067 ( .A1(n2060), .A2(n2061), .Y(n2045) );
  OR2X1_RVT U2068 ( .A1(n2007), .A2(n2062), .Y(n2061) );
  OR2X1_RVT U2069 ( .A1(n2063), .A2(n12907), .Y(n2062) );
  OR2X1_RVT U2070 ( .A1(n2064), .A2(n2065), .Y(n2060) );
  OR2X1_RVT U2071 ( .A1(n2066), .A2(n12594), .Y(n2065) );
  OR2X1_RVT U2072 ( .A1(n1942), .A2(n2067), .Y(n1935) );
  AND4X1_RVT U2073 ( .A1(n2068), .A2(n2069), .A3(n2070), .A4(n2071), .Y(n2042)
         );
  AND4X1_RVT U2074 ( .A1(n2072), .A2(n2073), .A3(n2074), .A4(n2075), .Y(n2071)
         );
  OR2X1_RVT U2075 ( .A1(n2076), .A2(n12608), .Y(n2075) );
  AND2X1_RVT U2076 ( .A1(n2078), .A2(n2079), .Y(n2076) );
  OR2X1_RVT U2077 ( .A1(n12577), .A2(n1957), .Y(n2079) );
  OR2X1_RVT U2078 ( .A1(n2080), .A2(n1959), .Y(n2074) );
  AND2X1_RVT U2079 ( .A1(n2081), .A2(n2082), .Y(n2080) );
  OR2X1_RVT U2080 ( .A1(n2083), .A2(n12906), .Y(n2073) );
  AND2X1_RVT U2081 ( .A1(n2084), .A2(n2085), .Y(n2083) );
  OR2X1_RVT U2082 ( .A1(n2086), .A2(n2035), .Y(n2085) );
  AND2X1_RVT U2083 ( .A1(n12608), .A2(n12592), .Y(n2086) );
  OR2X1_RVT U2084 ( .A1(n2087), .A2(n12578), .Y(n2072) );
  AND2X1_RVT U2085 ( .A1(n2089), .A2(n2090), .Y(n2087) );
  OR2X1_RVT U2086 ( .A1(n2091), .A2(n12584), .Y(n2070) );
  AND2X1_RVT U2087 ( .A1(n2092), .A2(n2093), .Y(n2091) );
  OR2X1_RVT U2088 ( .A1(n12592), .A2(n2094), .Y(n2093) );
  AND2X1_RVT U2089 ( .A1(n2095), .A2(n2096), .Y(n2092) );
  OR2X1_RVT U2090 ( .A1(n2097), .A2(n2098), .Y(n2095) );
  OR2X1_RVT U2091 ( .A1(n1942), .A2(n2013), .Y(n2098) );
  OR2X1_RVT U2092 ( .A1(n2099), .A2(n12903), .Y(n2069) );
  AND2X1_RVT U2093 ( .A1(n2100), .A2(n2101), .Y(n2099) );
  OR2X1_RVT U2094 ( .A1(n2102), .A2(n2103), .Y(n2068) );
  AND2X1_RVT U2095 ( .A1(n2104), .A2(n2105), .Y(n2102) );
  AND2X1_RVT U2096 ( .A1(n2106), .A2(n2107), .Y(n2104) );
  OR2X1_RVT U2097 ( .A1(n31), .A2(n2035), .Y(n2107) );
  OR2X1_RVT U2098 ( .A1(n12602), .A2(n2000), .Y(n2106) );
  AND4X1_RVT U2099 ( .A1(n2108), .A2(n2109), .A3(n2110), .A4(n2111), .Y(n2041)
         );
  AND4X1_RVT U2100 ( .A1(n2112), .A2(n2113), .A3(n2114), .A4(n2115), .Y(n2111)
         );
  OR2X1_RVT U2101 ( .A1(n2035), .A2(n2034), .Y(n2115) );
  OR2X1_RVT U2102 ( .A1(n1966), .A2(n2116), .Y(n2114) );
  OR2X1_RVT U2103 ( .A1(n1999), .A2(n2117), .Y(n2113) );
  OR2X1_RVT U2104 ( .A1(n1942), .A2(n2118), .Y(n2112) );
  AND2X1_RVT U2105 ( .A1(n2119), .A2(n2120), .Y(n2110) );
  OR2X1_RVT U2106 ( .A1(n12603), .A2(n2121), .Y(n2120) );
  OR2X1_RVT U2107 ( .A1(n12582), .A2(n2018), .Y(n2119) );
  OR2X1_RVT U2108 ( .A1(n2122), .A2(n1977), .Y(n2109) );
  AND4X1_RVT U2109 ( .A1(n2123), .A2(n2124), .A3(n2125), .A4(n2126), .Y(n2122)
         );
  OR2X1_RVT U2110 ( .A1(n2127), .A2(n1942), .Y(n2125) );
  OR2X1_RVT U2111 ( .A1(n12895), .A2(n2128), .Y(n2124) );
  OR2X1_RVT U2112 ( .A1(n2129), .A2(n12903), .Y(n2123) );
  AND2X1_RVT U2113 ( .A1(n2020), .A2(n2130), .Y(n2129) );
  OR2X1_RVT U2114 ( .A1(n2022), .A2(n2131), .Y(n2108) );
  AND4X1_RVT U2115 ( .A1(n2132), .A2(n2133), .A3(n2134), .A4(n2135), .Y(n2040)
         );
  AND4X1_RVT U2116 ( .A1(n2136), .A2(n2137), .A3(n2138), .A4(n2139), .Y(n2135)
         );
  OR2X1_RVT U2117 ( .A1(n12899), .A2(n2140), .Y(n2139) );
  OR2X1_RVT U2118 ( .A1(n12900), .A2(n2141), .Y(n2138) );
  OR2X1_RVT U2119 ( .A1(n12897), .A2(n2142), .Y(n2137) );
  OR2X1_RVT U2120 ( .A1(n12576), .A2(n2143), .Y(n2136) );
  OR2X1_RVT U2121 ( .A1(n2144), .A2(n12583), .Y(n2133) );
  AND4X1_RVT U2122 ( .A1(n2146), .A2(n2147), .A3(n2148), .A4(n2149), .Y(n2145)
         );
  AND4X1_RVT U2123 ( .A1(n2150), .A2(n2151), .A3(n2152), .A4(n2153), .Y(n2149)
         );
  AND4X1_RVT U2124 ( .A1(n2154), .A2(n1931), .A3(n2101), .A4(n2155), .Y(n2153)
         );
  OR2X1_RVT U2125 ( .A1(n2156), .A2(n12894), .Y(n1931) );
  AND2X1_RVT U2126 ( .A1(n2157), .A2(n2158), .Y(n2156) );
  OR2X1_RVT U2127 ( .A1(n1975), .A2(n2159), .Y(n2158) );
  OR2X1_RVT U2128 ( .A1(n2160), .A2(n2057), .Y(n2157) );
  OR2X1_RVT U2129 ( .A1(n2161), .A2(n2016), .Y(n2154) );
  AND2X1_RVT U2130 ( .A1(n2162), .A2(n2163), .Y(n2161) );
  OR2X1_RVT U2131 ( .A1(n12899), .A2(n2000), .Y(n2163) );
  OR2X1_RVT U2132 ( .A1(n2164), .A2(n1959), .Y(n2152) );
  AND2X1_RVT U2133 ( .A1(n2165), .A2(n2166), .Y(n2164) );
  OR2X1_RVT U2134 ( .A1(n2167), .A2(n12905), .Y(n2166) );
  AND2X1_RVT U2135 ( .A1(n2007), .A2(n2168), .Y(n2167) );
  OR2X1_RVT U2136 ( .A1(n2169), .A2(n12603), .Y(n2151) );
  AND2X1_RVT U2137 ( .A1(n2170), .A2(n2171), .Y(n2169) );
  OR2X1_RVT U2138 ( .A1(n2000), .A2(n1966), .Y(n2171) );
  OR2X1_RVT U2139 ( .A1(n2172), .A2(n12586), .Y(n2150) );
  AND2X1_RVT U2140 ( .A1(n2084), .A2(n2173), .Y(n2172) );
  OR2X1_RVT U2141 ( .A1(n2013), .A2(n2174), .Y(n2084) );
  AND4X1_RVT U2142 ( .A1(n2175), .A2(n2176), .A3(n2177), .A4(n2178), .Y(n2148)
         );
  OR2X1_RVT U2143 ( .A1(n2179), .A2(n12593), .Y(n2178) );
  AND2X1_RVT U2144 ( .A1(n2180), .A2(n2181), .Y(n2179) );
  OR2X1_RVT U2145 ( .A1(n2057), .A2(n1957), .Y(n2181) );
  AND2X1_RVT U2146 ( .A1(n2182), .A2(n2183), .Y(n2180) );
  OR2X1_RVT U2147 ( .A1(n2097), .A2(n2159), .Y(n2182) );
  AND2X1_RVT U2148 ( .A1(n2184), .A2(n2185), .Y(n2177) );
  OR2X1_RVT U2149 ( .A1(n2186), .A2(n2088), .Y(n2185) );
  AND2X1_RVT U2150 ( .A1(n2187), .A2(n1996), .Y(n2186) );
  OR2X1_RVT U2151 ( .A1(n1942), .A2(n2057), .Y(n1996) );
  OR2X1_RVT U2152 ( .A1(n2188), .A2(n31), .Y(n2184) );
  AND2X1_RVT U2153 ( .A1(n2189), .A2(n2190), .Y(n2188) );
  OR2X1_RVT U2154 ( .A1(n2191), .A2(n12595), .Y(n2190) );
  AND2X1_RVT U2155 ( .A1(n2192), .A2(n2193), .Y(n2191) );
  OR2X1_RVT U2156 ( .A1(n12590), .A2(n2007), .Y(n2193) );
  OR2X1_RVT U2157 ( .A1(n12909), .A2(n12592), .Y(n2192) );
  AND2X1_RVT U2158 ( .A1(n2058), .A2(n2168), .Y(n2189) );
  OR2X1_RVT U2159 ( .A1(n2088), .A2(n2194), .Y(n2058) );
  OR2X1_RVT U2160 ( .A1(n12904), .A2(n12900), .Y(n2194) );
  OR2X1_RVT U2161 ( .A1(n2195), .A2(n2077), .Y(n2176) );
  AND4X1_RVT U2162 ( .A1(n2036), .A2(n2196), .A3(n2197), .A4(n2198), .Y(n2195)
         );
  OR2X1_RVT U2163 ( .A1(n12594), .A2(n2057), .Y(n2198) );
  AND2X1_RVT U2164 ( .A1(n2199), .A2(n2200), .Y(n2197) );
  OR2X1_RVT U2165 ( .A1(n12909), .A2(n12603), .Y(n2196) );
  AND2X1_RVT U2166 ( .A1(n2201), .A2(n2202), .Y(n2036) );
  OR2X1_RVT U2167 ( .A1(n2203), .A2(n29), .Y(n2202) );
  OR2X1_RVT U2168 ( .A1(n2000), .A2(n12894), .Y(n2201) );
  AND2X1_RVT U2169 ( .A1(n2204), .A2(n2205), .Y(n2175) );
  OR2X1_RVT U2170 ( .A1(n2206), .A2(n12896), .Y(n2205) );
  AND2X1_RVT U2171 ( .A1(n2207), .A2(n2208), .Y(n2206) );
  OR2X1_RVT U2172 ( .A1(n2209), .A2(n12597), .Y(n2208) );
  AND2X1_RVT U2173 ( .A1(n2210), .A2(n2211), .Y(n2209) );
  AND2X1_RVT U2174 ( .A1(n2212), .A2(n2213), .Y(n2207) );
  OR2X1_RVT U2175 ( .A1(n2214), .A2(n12606), .Y(n2204) );
  AND4X1_RVT U2176 ( .A1(n2215), .A2(n2216), .A3(n2217), .A4(n2218), .Y(n2214)
         );
  OR2X1_RVT U2177 ( .A1(n12908), .A2(n2219), .Y(n2217) );
  OR2X1_RVT U2178 ( .A1(n29), .A2(n2014), .Y(n2216) );
  OR2X1_RVT U2179 ( .A1(n2103), .A2(n2057), .Y(n2215) );
  AND4X1_RVT U2180 ( .A1(n2220), .A2(n2221), .A3(n2222), .A4(n2223), .Y(n2147)
         );
  AND2X1_RVT U2181 ( .A1(n2224), .A2(n2067), .Y(n2223) );
  OR2X1_RVT U2182 ( .A1(n12581), .A2(n2033), .Y(n2067) );
  AND2X1_RVT U2183 ( .A1(n2225), .A2(n2226), .Y(n2224) );
  OR2X1_RVT U2184 ( .A1(n2227), .A2(n1982), .Y(n2226) );
  OR2X1_RVT U2185 ( .A1(n2034), .A2(n2094), .Y(n2225) );
  OR2X1_RVT U2186 ( .A1(n29), .A2(n2228), .Y(n2222) );
  OR2X1_RVT U2187 ( .A1(n12907), .A2(n2229), .Y(n2221) );
  OR2X1_RVT U2188 ( .A1(n2103), .A2(n2230), .Y(n2220) );
  AND4X1_RVT U2189 ( .A1(n2231), .A2(n2232), .A3(n2233), .A4(n2234), .Y(n2146)
         );
  AND2X1_RVT U2190 ( .A1(n2235), .A2(n2236), .Y(n2234) );
  OR2X1_RVT U2191 ( .A1(n12576), .A2(n2237), .Y(n2236) );
  AND2X1_RVT U2192 ( .A1(n2238), .A2(n2239), .Y(n2235) );
  OR2X1_RVT U2193 ( .A1(n1999), .A2(n2009), .Y(n2239) );
  OR2X1_RVT U2194 ( .A1(n12597), .A2(n2059), .Y(n2009) );
  OR2X1_RVT U2195 ( .A1(n12583), .A2(n2240), .Y(n2238) );
  OR2X1_RVT U2196 ( .A1(n1980), .A2(n1973), .Y(n2233) );
  OR2X1_RVT U2197 ( .A1(n2066), .A2(n2241), .Y(n1973) );
  OR2X1_RVT U2198 ( .A1(n12903), .A2(n2242), .Y(n2232) );
  OR2X1_RVT U2199 ( .A1(n12595), .A2(n2100), .Y(n2231) );
  OR2X1_RVT U2200 ( .A1(n12894), .A2(n2162), .Y(n2100) );
  AND4X1_RVT U2201 ( .A1(n2244), .A2(n2245), .A3(n2246), .A4(n2247), .Y(n2243)
         );
  AND4X1_RVT U2202 ( .A1(n2248), .A2(n2249), .A3(n2250), .A4(n2251), .Y(n2247)
         );
  OR2X1_RVT U2203 ( .A1(n39), .A2(n2252), .Y(n2251) );
  OR2X1_RVT U2204 ( .A1(n2253), .A2(n12608), .Y(n2252) );
  AND2X1_RVT U2205 ( .A1(n12597), .A2(n2019), .Y(n2253) );
  AND2X1_RVT U2206 ( .A1(n1934), .A2(n2254), .Y(n2250) );
  OR2X1_RVT U2207 ( .A1(n12586), .A2(n2255), .Y(n1934) );
  OR2X1_RVT U2208 ( .A1(n39), .A2(n2013), .Y(n2255) );
  OR2X1_RVT U2209 ( .A1(n2256), .A2(n1942), .Y(n2249) );
  AND2X1_RVT U2210 ( .A1(n2257), .A2(n2258), .Y(n2256) );
  AND2X1_RVT U2211 ( .A1(n2259), .A2(n2260), .Y(n2248) );
  OR2X1_RVT U2212 ( .A1(n2261), .A2(n2262), .Y(n2260) );
  AND2X1_RVT U2213 ( .A1(n2263), .A2(n2023), .Y(n2261) );
  OR2X1_RVT U2214 ( .A1(n2264), .A2(n2014), .Y(n2259) );
  AND2X1_RVT U2215 ( .A1(n2199), .A2(n2033), .Y(n2264) );
  OR2X1_RVT U2216 ( .A1(n12584), .A2(n2265), .Y(n2199) );
  OR2X1_RVT U2217 ( .A1(n12909), .A2(n12594), .Y(n2265) );
  AND4X1_RVT U2218 ( .A1(n2266), .A2(n2267), .A3(n2268), .A4(n2269), .Y(n2246)
         );
  OR2X1_RVT U2219 ( .A1(n2270), .A2(n12899), .Y(n2269) );
  AND2X1_RVT U2220 ( .A1(n2082), .A2(n2271), .Y(n2270) );
  OR2X1_RVT U2221 ( .A1(n12907), .A2(n2127), .Y(n2082) );
  AND2X1_RVT U2222 ( .A1(n2272), .A2(n2273), .Y(n2268) );
  OR2X1_RVT U2223 ( .A1(n2274), .A2(n12897), .Y(n2273) );
  AND2X1_RVT U2224 ( .A1(n2275), .A2(n2276), .Y(n2274) );
  OR2X1_RVT U2225 ( .A1(n1977), .A2(n2219), .Y(n2276) );
  OR2X1_RVT U2226 ( .A1(n2277), .A2(n12895), .Y(n2272) );
  AND2X1_RVT U2227 ( .A1(n2278), .A2(n2279), .Y(n2277) );
  OR2X1_RVT U2228 ( .A1(n2280), .A2(n12597), .Y(n2267) );
  AND2X1_RVT U2229 ( .A1(n2281), .A2(n2282), .Y(n2280) );
  AND2X1_RVT U2230 ( .A1(n2283), .A2(n2284), .Y(n2281) );
  AND2X1_RVT U2231 ( .A1(n2285), .A2(n2286), .Y(n2266) );
  OR2X1_RVT U2232 ( .A1(n2287), .A2(n2203), .Y(n2286) );
  AND2X1_RVT U2233 ( .A1(n2288), .A2(n2034), .Y(n2287) );
  AND2X1_RVT U2234 ( .A1(n2289), .A2(n2290), .Y(n2288) );
  OR2X1_RVT U2235 ( .A1(n2291), .A2(n12600), .Y(n2285) );
  AND2X1_RVT U2236 ( .A1(n2292), .A2(n2293), .Y(n2291) );
  OR2X1_RVT U2237 ( .A1(n12906), .A2(n12602), .Y(n2293) );
  AND2X1_RVT U2238 ( .A1(n2023), .A2(n2294), .Y(n2292) );
  AND4X1_RVT U2239 ( .A1(n2295), .A2(n2296), .A3(n2297), .A4(n2298), .Y(n2245)
         );
  AND2X1_RVT U2240 ( .A1(n2299), .A2(n2300), .Y(n2298) );
  OR2X1_RVT U2241 ( .A1(n2016), .A2(n2090), .Y(n2300) );
  OR2X1_RVT U2242 ( .A1(n12901), .A2(n2023), .Y(n2090) );
  AND2X1_RVT U2243 ( .A1(n2301), .A2(n2302), .Y(n2299) );
  OR2X1_RVT U2244 ( .A1(n2168), .A2(n1982), .Y(n2302) );
  OR2X1_RVT U2245 ( .A1(n12908), .A2(n12593), .Y(n1982) );
  OR2X1_RVT U2246 ( .A1(n2066), .A2(n2116), .Y(n2301) );
  OR2X1_RVT U2247 ( .A1(n12896), .A2(n2303), .Y(n2116) );
  OR2X1_RVT U2248 ( .A1(n2304), .A2(n12576), .Y(n2297) );
  AND4X1_RVT U2249 ( .A1(n2305), .A2(n2306), .A3(n2307), .A4(n2308), .Y(n2304)
         );
  OR2X1_RVT U2250 ( .A1(n2241), .A2(n2014), .Y(n2307) );
  OR2X1_RVT U2251 ( .A1(n2309), .A2(n2011), .Y(n2306) );
  OR2X1_RVT U2252 ( .A1(n12905), .A2(n1966), .Y(n2305) );
  OR2X1_RVT U2253 ( .A1(n2310), .A2(n12577), .Y(n2296) );
  AND2X1_RVT U2254 ( .A1(n2311), .A2(n2312), .Y(n2310) );
  OR2X1_RVT U2255 ( .A1(n2241), .A2(n1966), .Y(n2312) );
  AND2X1_RVT U2256 ( .A1(n2313), .A2(n2242), .Y(n2311) );
  OR2X1_RVT U2257 ( .A1(n2014), .A2(n2314), .Y(n2242) );
  OR2X1_RVT U2258 ( .A1(n12896), .A2(n12908), .Y(n2314) );
  OR2X1_RVT U2259 ( .A1(n2315), .A2(n12584), .Y(n2295) );
  AND4X1_RVT U2260 ( .A1(n2316), .A2(n2229), .A3(n2038), .A4(n2010), .Y(n2315)
         );
  OR2X1_RVT U2261 ( .A1(n2035), .A2(n2317), .Y(n2010) );
  OR2X1_RVT U2262 ( .A1(n12898), .A2(n1972), .Y(n2317) );
  OR2X1_RVT U2263 ( .A1(n2097), .A2(n2131), .Y(n2038) );
  OR2X1_RVT U2264 ( .A1(n2016), .A2(n2318), .Y(n2229) );
  OR2X1_RVT U2265 ( .A1(n12608), .A2(n12577), .Y(n2318) );
  OR2X1_RVT U2266 ( .A1(n1975), .A2(n2319), .Y(n2316) );
  OR2X1_RVT U2267 ( .A1(n2320), .A2(n12582), .Y(n2319) );
  AND4X1_RVT U2268 ( .A1(n2321), .A2(n2322), .A3(n2323), .A4(n2324), .Y(n2244)
         );
  AND2X1_RVT U2269 ( .A1(n2325), .A2(n2326), .Y(n2324) );
  AND2X1_RVT U2270 ( .A1(n2327), .A2(n2328), .Y(n2325) );
  OR2X1_RVT U2271 ( .A1(n2007), .A2(n2282), .Y(n2328) );
  OR2X1_RVT U2272 ( .A1(n2019), .A2(n2329), .Y(n2282) );
  OR2X1_RVT U2273 ( .A1(n12897), .A2(n12899), .Y(n2329) );
  OR2X1_RVT U2274 ( .A1(n12904), .A2(n2330), .Y(n2327) );
  OR2X1_RVT U2275 ( .A1(n12593), .A2(n2331), .Y(n2323) );
  OR2X1_RVT U2276 ( .A1(n12907), .A2(n2332), .Y(n2322) );
  OR2X1_RVT U2277 ( .A1(n2019), .A2(n2333), .Y(n2321) );
  AND4X1_RVT U2278 ( .A1(n2335), .A2(n2336), .A3(n2337), .A4(n2338), .Y(n2334)
         );
  AND4X1_RVT U2279 ( .A1(n2339), .A2(n2340), .A3(n2341), .A4(n2342), .Y(n2338)
         );
  AND4X1_RVT U2280 ( .A1(n2343), .A2(n2344), .A3(n1936), .A4(n2345), .Y(n2342)
         );
  OR2X1_RVT U2281 ( .A1(n2077), .A2(n2346), .Y(n1936) );
  OR2X1_RVT U2282 ( .A1(n2168), .A2(n31), .Y(n2346) );
  OR2X1_RVT U2283 ( .A1(n1940), .A2(n2347), .Y(n2344) );
  OR2X1_RVT U2284 ( .A1(n12902), .A2(n12905), .Y(n2347) );
  OR2X1_RVT U2285 ( .A1(n2203), .A2(n2348), .Y(n2343) );
  OR2X1_RVT U2286 ( .A1(n2349), .A2(n1977), .Y(n2348) );
  AND2X1_RVT U2287 ( .A1(n12597), .A2(n2077), .Y(n2349) );
  OR2X1_RVT U2288 ( .A1(n2350), .A2(n12603), .Y(n2341) );
  AND2X1_RVT U2289 ( .A1(n2218), .A2(n2290), .Y(n2350) );
  OR2X1_RVT U2290 ( .A1(n31), .A2(n2351), .Y(n2290) );
  OR2X1_RVT U2291 ( .A1(n12576), .A2(n12901), .Y(n2351) );
  OR2X1_RVT U2292 ( .A1(n2007), .A2(n2352), .Y(n2218) );
  OR2X1_RVT U2293 ( .A1(n12899), .A2(n1999), .Y(n2352) );
  OR2X1_RVT U2294 ( .A1(n2353), .A2(n1957), .Y(n2340) );
  AND2X1_RVT U2295 ( .A1(n2354), .A2(n2162), .Y(n2353) );
  OR2X1_RVT U2296 ( .A1(n2063), .A2(n2057), .Y(n2339) );
  AND4X1_RVT U2297 ( .A1(n2355), .A2(n2356), .A3(n2357), .A4(n2358), .Y(n2337)
         );
  AND2X1_RVT U2298 ( .A1(n2359), .A2(n2360), .Y(n2358) );
  OR2X1_RVT U2299 ( .A1(n2361), .A2(n12597), .Y(n2360) );
  AND2X1_RVT U2300 ( .A1(n2362), .A2(n2030), .Y(n2361) );
  AND2X1_RVT U2301 ( .A1(n2363), .A2(n2364), .Y(n2359) );
  OR2X1_RVT U2302 ( .A1(n2365), .A2(n2013), .Y(n2364) );
  AND2X1_RVT U2303 ( .A1(n1984), .A2(n1956), .Y(n2365) );
  OR2X1_RVT U2304 ( .A1(n12907), .A2(n2055), .Y(n1984) );
  OR2X1_RVT U2305 ( .A1(n2366), .A2(n2066), .Y(n2363) );
  AND2X1_RVT U2306 ( .A1(n2258), .A2(n2367), .Y(n2366) );
  OR2X1_RVT U2307 ( .A1(n12908), .A2(n2094), .Y(n2258) );
  OR2X1_RVT U2308 ( .A1(n2368), .A2(n12899), .Y(n2357) );
  AND2X1_RVT U2309 ( .A1(n1961), .A2(n2369), .Y(n2368) );
  OR2X1_RVT U2310 ( .A1(n2097), .A2(n2021), .Y(n2369) );
  OR2X1_RVT U2311 ( .A1(n2000), .A2(n2203), .Y(n1961) );
  OR2X1_RVT U2312 ( .A1(n2370), .A2(n29), .Y(n2356) );
  AND2X1_RVT U2313 ( .A1(n2011), .A2(n2371), .Y(n2370) );
  OR2X1_RVT U2314 ( .A1(n2372), .A2(n12581), .Y(n2371) );
  AND2X1_RVT U2315 ( .A1(n2373), .A2(n2374), .Y(n2372) );
  OR2X1_RVT U2316 ( .A1(n12900), .A2(n1994), .Y(n2374) );
  OR2X1_RVT U2317 ( .A1(n12608), .A2(n2097), .Y(n2011) );
  OR2X1_RVT U2318 ( .A1(n2375), .A2(n2081), .Y(n2355) );
  AND2X1_RVT U2319 ( .A1(n2014), .A2(n2059), .Y(n2375) );
  OR2X1_RVT U2320 ( .A1(n12896), .A2(n1942), .Y(n2059) );
  AND4X1_RVT U2321 ( .A1(n2376), .A2(n2377), .A3(n2378), .A4(n2379), .Y(n2336)
         );
  AND4X1_RVT U2322 ( .A1(n2380), .A2(n2381), .A3(n2382), .A4(n2383), .Y(n2379)
         );
  OR2X1_RVT U2323 ( .A1(n2384), .A2(n12907), .Y(n2383) );
  AND2X1_RVT U2324 ( .A1(n2117), .A2(n2385), .Y(n2384) );
  OR2X1_RVT U2325 ( .A1(n12605), .A2(n1966), .Y(n2385) );
  OR2X1_RVT U2326 ( .A1(n2386), .A2(n1959), .Y(n2382) );
  AND2X1_RVT U2327 ( .A1(n2387), .A2(n2388), .Y(n2386) );
  OR2X1_RVT U2328 ( .A1(n2389), .A2(n1994), .Y(n2388) );
  AND2X1_RVT U2329 ( .A1(n2019), .A2(n2007), .Y(n2389) );
  AND2X1_RVT U2330 ( .A1(n2021), .A2(n2263), .Y(n2387) );
  OR2X1_RVT U2331 ( .A1(n12606), .A2(n2159), .Y(n2263) );
  OR2X1_RVT U2332 ( .A1(n2390), .A2(n12595), .Y(n2381) );
  AND2X1_RVT U2333 ( .A1(n2391), .A2(n2392), .Y(n2390) );
  OR2X1_RVT U2334 ( .A1(n2007), .A2(n2393), .Y(n2392) );
  AND2X1_RVT U2335 ( .A1(n2089), .A2(n2283), .Y(n2391) );
  OR2X1_RVT U2336 ( .A1(n1999), .A2(n2174), .Y(n2283) );
  OR2X1_RVT U2337 ( .A1(n1972), .A2(n2394), .Y(n2089) );
  OR2X1_RVT U2338 ( .A1(n2395), .A2(n1942), .Y(n2380) );
  AND4X1_RVT U2339 ( .A1(n2396), .A2(n2397), .A3(n2398), .A4(n2331), .Y(n2395)
         );
  OR2X1_RVT U2340 ( .A1(n2035), .A2(n2399), .Y(n2331) );
  OR2X1_RVT U2341 ( .A1(n12576), .A2(n1999), .Y(n2399) );
  OR2X1_RVT U2342 ( .A1(n12904), .A2(n2241), .Y(n2397) );
  OR2X1_RVT U2343 ( .A1(n2000), .A2(n2097), .Y(n2396) );
  OR2X1_RVT U2344 ( .A1(n2168), .A2(n2210), .Y(n2378) );
  OR2X1_RVT U2345 ( .A1(n2400), .A2(n12579), .Y(n2377) );
  AND4X1_RVT U2346 ( .A1(n2401), .A2(n2402), .A3(n2044), .A4(n2142), .Y(n2400)
         );
  OR2X1_RVT U2347 ( .A1(n1966), .A2(n2131), .Y(n2142) );
  OR2X1_RVT U2348 ( .A1(n12904), .A2(n29), .Y(n2131) );
  OR2X1_RVT U2349 ( .A1(n1959), .A2(n2023), .Y(n2044) );
  OR2X1_RVT U2350 ( .A1(n12896), .A2(n2394), .Y(n2376) );
  AND4X1_RVT U2351 ( .A1(n2403), .A2(n2404), .A3(n2405), .A4(n2406), .Y(n2335)
         );
  OR2X1_RVT U2352 ( .A1(n12584), .A2(n2407), .Y(n2406) );
  AND2X1_RVT U2353 ( .A1(n2408), .A2(n2409), .Y(n2405) );
  OR2X1_RVT U2354 ( .A1(n12605), .A2(n2162), .Y(n2409) );
  OR2X1_RVT U2355 ( .A1(n1949), .A2(n2023), .Y(n2408) );
  OR2X1_RVT U2356 ( .A1(n31), .A2(n1980), .Y(n2023) );
  OR2X1_RVT U2357 ( .A1(n12608), .A2(n2141), .Y(n2404) );
  OR2X1_RVT U2358 ( .A1(n2016), .A2(n2410), .Y(n2141) );
  AND2X1_RVT U2359 ( .A1(n2411), .A2(n2412), .Y(n2403) );
  OR2X1_RVT U2360 ( .A1(n12577), .A2(n2413), .Y(n2412) );
  OR2X1_RVT U2361 ( .A1(n2019), .A2(n1968), .Y(n2411) );
  OR2X1_RVT U2362 ( .A1(n1942), .A2(n2227), .Y(n1968) );
  AND4X1_RVT U2363 ( .A1(n2415), .A2(n2416), .A3(n2417), .A4(n2418), .Y(n2414)
         );
  AND4X1_RVT U2364 ( .A1(n2419), .A2(n2420), .A3(n2421), .A4(n2422), .Y(n2418)
         );
  AND4X1_RVT U2365 ( .A1(n2155), .A2(n2345), .A3(n2423), .A4(n2424), .Y(n2422)
         );
  OR2X1_RVT U2366 ( .A1(n2425), .A2(n2426), .Y(n2345) );
  OR2X1_RVT U2367 ( .A1(n1940), .A2(n2210), .Y(n2155) );
  OR2X1_RVT U2368 ( .A1(n12905), .A2(n12593), .Y(n2210) );
  AND4X1_RVT U2369 ( .A1(n2413), .A2(n2279), .A3(n2402), .A4(n1937), .Y(n2421)
         );
  OR2X1_RVT U2370 ( .A1(n2427), .A2(n2127), .Y(n1937) );
  OR2X1_RVT U2371 ( .A1(n1942), .A2(n2428), .Y(n2402) );
  OR2X1_RVT U2372 ( .A1(n1975), .A2(n29), .Y(n2279) );
  OR2X1_RVT U2373 ( .A1(n1966), .A2(n2429), .Y(n2413) );
  OR2X1_RVT U2374 ( .A1(n12583), .A2(n12603), .Y(n2429) );
  AND4X1_RVT U2375 ( .A1(n2430), .A2(n2431), .A3(n2432), .A4(n2433), .Y(n2420)
         );
  OR2X1_RVT U2376 ( .A1(n2219), .A2(n2434), .Y(n2433) );
  OR2X1_RVT U2377 ( .A1(n12603), .A2(n1999), .Y(n2434) );
  OR2X1_RVT U2378 ( .A1(n2128), .A2(n2435), .Y(n2432) );
  OR2X1_RVT U2379 ( .A1(n12906), .A2(n2016), .Y(n2435) );
  OR2X1_RVT U2380 ( .A1(n2354), .A2(n2436), .Y(n2431) );
  OR2X1_RVT U2381 ( .A1(n2437), .A2(n2013), .Y(n2436) );
  OR2X1_RVT U2382 ( .A1(n12600), .A2(n2438), .Y(n2430) );
  OR2X1_RVT U2383 ( .A1(n2439), .A2(n12583), .Y(n2438) );
  AND2X1_RVT U2384 ( .A1(n2227), .A2(n2440), .Y(n2439) );
  AND2X1_RVT U2385 ( .A1(n2441), .A2(n2442), .Y(n2419) );
  OR2X1_RVT U2386 ( .A1(n2443), .A2(n1994), .Y(n2442) );
  AND2X1_RVT U2387 ( .A1(n2444), .A2(n2445), .Y(n2443) );
  OR2X1_RVT U2388 ( .A1(n12582), .A2(n2187), .Y(n2445) );
  OR2X1_RVT U2389 ( .A1(n12586), .A2(n2262), .Y(n2444) );
  AND2X1_RVT U2390 ( .A1(n2446), .A2(n2447), .Y(n2441) );
  OR2X1_RVT U2391 ( .A1(n2448), .A2(n2033), .Y(n2447) );
  AND2X1_RVT U2392 ( .A1(n2449), .A2(n2450), .Y(n2448) );
  OR2X1_RVT U2393 ( .A1(n12589), .A2(n39), .Y(n2450) );
  NAND2X1_RVT U2394 ( .A1(n2016), .A2(n12898), .Y(n2449) );
  OR2X1_RVT U2395 ( .A1(n2451), .A2(n31), .Y(n2446) );
  AND2X1_RVT U2396 ( .A1(n2240), .A2(n2117), .Y(n2451) );
  OR2X1_RVT U2397 ( .A1(n1966), .A2(n2452), .Y(n2117) );
  OR2X1_RVT U2398 ( .A1(n12909), .A2(n12578), .Y(n2452) );
  AND4X1_RVT U2399 ( .A1(n2134), .A2(n2453), .A3(n2326), .A4(n2454), .Y(n2417)
         );
  AND4X1_RVT U2400 ( .A1(n2455), .A2(n2456), .A3(n2457), .A4(n2458), .Y(n2454)
         );
  OR2X1_RVT U2401 ( .A1(n2097), .A2(n2018), .Y(n2458) );
  OR2X1_RVT U2402 ( .A1(n2035), .A2(n2064), .Y(n2457) );
  OR2X1_RVT U2403 ( .A1(n12897), .A2(n2289), .Y(n2456) );
  OR2X1_RVT U2404 ( .A1(n2013), .A2(n1995), .Y(n2289) );
  OR2X1_RVT U2405 ( .A1(n12905), .A2(n2077), .Y(n1995) );
  OR2X1_RVT U2406 ( .A1(n12592), .A2(n2118), .Y(n2455) );
  OR2X1_RVT U2407 ( .A1(n1999), .A2(n2227), .Y(n2118) );
  OR2X1_RVT U2408 ( .A1(n12576), .A2(n2203), .Y(n2227) );
  AND2X1_RVT U2409 ( .A1(n2459), .A2(n2460), .Y(n2326) );
  OR2X1_RVT U2410 ( .A1(n2461), .A2(n2066), .Y(n2460) );
  OR2X1_RVT U2411 ( .A1(n12602), .A2(n31), .Y(n2461) );
  OR2X1_RVT U2412 ( .A1(n2462), .A2(n1949), .Y(n2459) );
  OR2X1_RVT U2413 ( .A1(n12896), .A2(n2066), .Y(n1949) );
  OR2X1_RVT U2414 ( .A1(n1963), .A2(n2013), .Y(n2462) );
  OR2X1_RVT U2415 ( .A1(n12584), .A2(n2332), .Y(n2453) );
  AND2X1_RVT U2416 ( .A1(n2463), .A2(n2464), .Y(n2134) );
  OR2X1_RVT U2417 ( .A1(n2017), .A2(n2055), .Y(n2464) );
  OR2X1_RVT U2418 ( .A1(n2465), .A2(n2466), .Y(n2463) );
  AND4X1_RVT U2419 ( .A1(n2467), .A2(n2468), .A3(n2469), .A4(n2470), .Y(n2416)
         );
  OR2X1_RVT U2420 ( .A1(n2471), .A2(n2203), .Y(n2470) );
  AND2X1_RVT U2421 ( .A1(n2472), .A2(n2212), .Y(n2471) );
  OR2X1_RVT U2422 ( .A1(n12590), .A2(n2428), .Y(n2212) );
  OR2X1_RVT U2423 ( .A1(n2473), .A2(n12902), .Y(n2469) );
  AND2X1_RVT U2424 ( .A1(n2140), .A2(n2105), .Y(n2473) );
  OR2X1_RVT U2425 ( .A1(n12896), .A2(n2081), .Y(n2105) );
  OR2X1_RVT U2426 ( .A1(n2474), .A2(n2160), .Y(n2468) );
  AND2X1_RVT U2427 ( .A1(n2475), .A2(n2476), .Y(n2474) );
  OR2X1_RVT U2428 ( .A1(n12579), .A2(n2019), .Y(n2476) );
  AND2X1_RVT U2429 ( .A1(n2477), .A2(n2057), .Y(n2475) );
  OR2X1_RVT U2430 ( .A1(n29), .A2(n2016), .Y(n2477) );
  OR2X1_RVT U2431 ( .A1(n2478), .A2(n1957), .Y(n2467) );
  AND2X1_RVT U2432 ( .A1(n2479), .A2(n2480), .Y(n2478) );
  NAND2X1_RVT U2433 ( .A1(n1942), .A2(n2320), .Y(n2480) );
  AND2X1_RVT U2434 ( .A1(n2481), .A2(n2170), .Y(n2479) );
  OR2X1_RVT U2435 ( .A1(n2103), .A2(n2428), .Y(n2170) );
  OR2X1_RVT U2436 ( .A1(n12599), .A2(n2482), .Y(n2481) );
  AND4X1_RVT U2437 ( .A1(n2483), .A2(n2484), .A3(n2485), .A4(n2486), .Y(n2415)
         );
  OR2X1_RVT U2438 ( .A1(n2487), .A2(n1980), .Y(n2486) );
  AND2X1_RVT U2439 ( .A1(n2488), .A2(n2121), .Y(n2487) );
  AND2X1_RVT U2440 ( .A1(n2489), .A2(n2143), .Y(n2488) );
  OR2X1_RVT U2441 ( .A1(n31), .A2(n2466), .Y(n2143) );
  OR2X1_RVT U2442 ( .A1(n12578), .A2(n2077), .Y(n2466) );
  OR2X1_RVT U2443 ( .A1(n2490), .A2(n12595), .Y(n2485) );
  AND2X1_RVT U2444 ( .A1(n2491), .A2(n2492), .Y(n2490) );
  OR2X1_RVT U2445 ( .A1(n2493), .A2(n12894), .Y(n2492) );
  AND2X1_RVT U2446 ( .A1(n2494), .A2(n2495), .Y(n2493) );
  OR2X1_RVT U2447 ( .A1(n12577), .A2(n2354), .Y(n2495) );
  OR2X1_RVT U2448 ( .A1(n12901), .A2(n2000), .Y(n2494) );
  AND2X1_RVT U2449 ( .A1(n2496), .A2(n2497), .Y(n2491) );
  OR2X1_RVT U2450 ( .A1(n1966), .A2(n2498), .Y(n2496) );
  OR2X1_RVT U2451 ( .A1(n2499), .A2(n2000), .Y(n2484) );
  AND4X1_RVT U2452 ( .A1(n2500), .A2(n2501), .A3(n2502), .A4(n1966), .Y(n2499)
         );
  OR2X1_RVT U2453 ( .A1(n12902), .A2(n2016), .Y(n2502) );
  OR2X1_RVT U2454 ( .A1(n12589), .A2(n2035), .Y(n2501) );
  OR2X1_RVT U2455 ( .A1(n2088), .A2(n2066), .Y(n2500) );
  OR2X1_RVT U2456 ( .A1(n2503), .A2(n1942), .Y(n2483) );
  AND4X1_RVT U2457 ( .A1(n2367), .A2(n2504), .A3(n2165), .A4(n2081), .Y(n2503)
         );
  OR2X1_RVT U2458 ( .A1(n2035), .A2(n2498), .Y(n2165) );
  OR2X1_RVT U2459 ( .A1(n2203), .A2(n2410), .Y(n2504) );
  OR2X1_RVT U2460 ( .A1(n12583), .A2(n2168), .Y(n2367) );
  AND4X1_RVT U2461 ( .A1(n2506), .A2(n2507), .A3(n2508), .A4(n2509), .Y(n2505)
         );
  AND4X1_RVT U2462 ( .A1(n2018), .A2(n2254), .A3(n2510), .A4(n2511), .Y(n2509)
         );
  AND4X1_RVT U2463 ( .A1(n2333), .A2(n2278), .A3(n2423), .A4(n2424), .Y(n2511)
         );
  OR2X1_RVT U2464 ( .A1(n2426), .A2(n1939), .Y(n2424) );
  OR2X1_RVT U2465 ( .A1(n12900), .A2(n2057), .Y(n1939) );
  OR2X1_RVT U2466 ( .A1(n1956), .A2(n2465), .Y(n2423) );
  OR2X1_RVT U2467 ( .A1(n12905), .A2(n12597), .Y(n2465) );
  OR2X1_RVT U2468 ( .A1(n12894), .A2(n2077), .Y(n1956) );
  OR2X1_RVT U2469 ( .A1(n12906), .A2(n1975), .Y(n2278) );
  OR2X1_RVT U2470 ( .A1(n12606), .A2(n12590), .Y(n1975) );
  OR2X1_RVT U2471 ( .A1(n2097), .A2(n2512), .Y(n2333) );
  OR2X1_RVT U2472 ( .A1(n12597), .A2(n2001), .Y(n2512) );
  OR2X1_RVT U2473 ( .A1(n1999), .A2(n2513), .Y(n2510) );
  OR2X1_RVT U2474 ( .A1(n2127), .A2(n12588), .Y(n2513) );
  OR2X1_RVT U2475 ( .A1(n2066), .A2(n2514), .Y(n2254) );
  OR2X1_RVT U2476 ( .A1(n2000), .A2(n12595), .Y(n2514) );
  OR2X1_RVT U2477 ( .A1(n12898), .A2(n2425), .Y(n2018) );
  OR2X1_RVT U2478 ( .A1(n12590), .A2(n2017), .Y(n2425) );
  AND4X1_RVT U2479 ( .A1(n2515), .A2(n2516), .A3(n2517), .A4(n2518), .Y(n2508)
         );
  AND4X1_RVT U2480 ( .A1(n2519), .A2(n2520), .A3(n2521), .A4(n2522), .Y(n2518)
         );
  OR2X1_RVT U2481 ( .A1(n2033), .A2(n2523), .Y(n2522) );
  OR2X1_RVT U2482 ( .A1(n12579), .A2(n2103), .Y(n2523) );
  OR2X1_RVT U2483 ( .A1(n2016), .A2(n2524), .Y(n2521) );
  OR2X1_RVT U2484 ( .A1(n2525), .A2(n1980), .Y(n2524) );
  AND2X1_RVT U2485 ( .A1(n1959), .A2(n2019), .Y(n2525) );
  OR2X1_RVT U2486 ( .A1(n2526), .A2(n2527), .Y(n2520) );
  AND2X1_RVT U2487 ( .A1(n2174), .A2(n2130), .Y(n2526) );
  OR2X1_RVT U2488 ( .A1(n12899), .A2(n39), .Y(n2130) );
  OR2X1_RVT U2489 ( .A1(n12895), .A2(n12600), .Y(n2174) );
  OR2X1_RVT U2490 ( .A1(n2528), .A2(n2014), .Y(n2519) );
  AND2X1_RVT U2491 ( .A1(n2410), .A2(n2529), .Y(n2528) );
  OR2X1_RVT U2492 ( .A1(n12897), .A2(n31), .Y(n2529) );
  OR2X1_RVT U2493 ( .A1(n2530), .A2(n12602), .Y(n2517) );
  AND2X1_RVT U2494 ( .A1(n2401), .A2(n2531), .Y(n2530) );
  OR2X1_RVT U2495 ( .A1(n2007), .A2(n2354), .Y(n2531) );
  OR2X1_RVT U2496 ( .A1(n12583), .A2(n2219), .Y(n2401) );
  OR2X1_RVT U2497 ( .A1(n12901), .A2(n2007), .Y(n2219) );
  OR2X1_RVT U2498 ( .A1(n2532), .A2(n2168), .Y(n2516) );
  AND2X1_RVT U2499 ( .A1(n2121), .A2(n2393), .Y(n2532) );
  OR2X1_RVT U2500 ( .A1(n1977), .A2(n2066), .Y(n2121) );
  OR2X1_RVT U2501 ( .A1(n2533), .A2(n2057), .Y(n2515) );
  AND2X1_RVT U2502 ( .A1(n2020), .A2(n2022), .Y(n2533) );
  AND4X1_RVT U2503 ( .A1(n2534), .A2(n2535), .A3(n2536), .A4(n2537), .Y(n2507)
         );
  AND4X1_RVT U2504 ( .A1(n2538), .A2(n2539), .A3(n2540), .A4(n2541), .Y(n2537)
         );
  OR2X1_RVT U2505 ( .A1(n2542), .A2(n12586), .Y(n2541) );
  AND2X1_RVT U2506 ( .A1(n1948), .A2(n2240), .Y(n2542) );
  OR2X1_RVT U2507 ( .A1(n2097), .A2(n2128), .Y(n2240) );
  OR2X1_RVT U2508 ( .A1(n12589), .A2(n1980), .Y(n2128) );
  OR2X1_RVT U2509 ( .A1(n12593), .A2(n2543), .Y(n1948) );
  OR2X1_RVT U2510 ( .A1(n12576), .A2(n12582), .Y(n2543) );
  OR2X1_RVT U2511 ( .A1(n2544), .A2(n12600), .Y(n2540) );
  AND2X1_RVT U2512 ( .A1(n2257), .A2(n2545), .Y(n2544) );
  OR2X1_RVT U2513 ( .A1(n12605), .A2(n29), .Y(n2545) );
  OR2X1_RVT U2514 ( .A1(n12603), .A2(n2064), .Y(n2257) );
  OR2X1_RVT U2515 ( .A1(n2546), .A2(n12581), .Y(n2539) );
  AND2X1_RVT U2516 ( .A1(n2275), .A2(n2547), .Y(n2546) );
  OR2X1_RVT U2517 ( .A1(n12606), .A2(n2000), .Y(n2547) );
  OR2X1_RVT U2518 ( .A1(n1942), .A2(n2548), .Y(n2275) );
  OR2X1_RVT U2519 ( .A1(n2549), .A2(n2001), .Y(n2538) );
  AND2X1_RVT U2520 ( .A1(n2550), .A2(n2551), .Y(n2549) );
  OR2X1_RVT U2521 ( .A1(n2057), .A2(n12603), .Y(n2551) );
  AND2X1_RVT U2522 ( .A1(n2552), .A2(n2033), .Y(n2550) );
  OR2X1_RVT U2523 ( .A1(n2019), .A2(n1980), .Y(n2033) );
  OR2X1_RVT U2524 ( .A1(n12578), .A2(n2064), .Y(n2552) );
  OR2X1_RVT U2525 ( .A1(n12909), .A2(n2019), .Y(n2064) );
  OR2X1_RVT U2526 ( .A1(n2553), .A2(n2077), .Y(n2536) );
  AND4X1_RVT U2527 ( .A1(n2554), .A2(n2555), .A3(n2230), .A4(n2140), .Y(n2553)
         );
  OR2X1_RVT U2528 ( .A1(n2203), .A2(n2303), .Y(n2140) );
  OR2X1_RVT U2529 ( .A1(n2035), .A2(n2482), .Y(n2230) );
  OR2X1_RVT U2530 ( .A1(n12584), .A2(n12577), .Y(n2482) );
  OR2X1_RVT U2531 ( .A1(n31), .A2(n1957), .Y(n2555) );
  OR2X1_RVT U2532 ( .A1(n29), .A2(n12603), .Y(n2554) );
  OR2X1_RVT U2533 ( .A1(n2556), .A2(n2013), .Y(n2535) );
  AND2X1_RVT U2534 ( .A1(n2557), .A2(n2034), .Y(n2556) );
  AND2X1_RVT U2535 ( .A1(n2489), .A2(n2284), .Y(n2557) );
  OR2X1_RVT U2536 ( .A1(n2558), .A2(n12906), .Y(n2284) );
  AND2X1_RVT U2537 ( .A1(n2055), .A2(n2559), .Y(n2558) );
  OR2X1_RVT U2538 ( .A1(n12581), .A2(n1942), .Y(n2559) );
  OR2X1_RVT U2539 ( .A1(n2103), .A2(n2241), .Y(n2489) );
  OR2X1_RVT U2540 ( .A1(n2088), .A2(n1977), .Y(n2241) );
  OR2X1_RVT U2541 ( .A1(n2560), .A2(n2081), .Y(n2534) );
  AND2X1_RVT U2542 ( .A1(n2561), .A2(n12589), .Y(n2560) );
  AND2X1_RVT U2543 ( .A1(n2562), .A2(n2262), .Y(n2561) );
  OR2X1_RVT U2544 ( .A1(n2103), .A2(n2203), .Y(n2562) );
  AND4X1_RVT U2545 ( .A1(n2563), .A2(n2564), .A3(n2565), .A4(n2566), .Y(n2506)
         );
  AND2X1_RVT U2546 ( .A1(n2567), .A2(n2568), .Y(n2566) );
  OR2X1_RVT U2547 ( .A1(n12902), .A2(n2183), .Y(n2568) );
  OR2X1_RVT U2548 ( .A1(n12597), .A2(n2569), .Y(n2183) );
  OR2X1_RVT U2549 ( .A1(n1999), .A2(n2088), .Y(n2569) );
  AND2X1_RVT U2550 ( .A1(n2570), .A2(n2571), .Y(n2567) );
  OR2X1_RVT U2551 ( .A1(n1972), .A2(n1983), .Y(n2571) );
  OR2X1_RVT U2552 ( .A1(n2016), .A2(n2211), .Y(n1983) );
  OR2X1_RVT U2553 ( .A1(n12898), .A2(n1977), .Y(n2211) );
  OR2X1_RVT U2554 ( .A1(n2019), .A2(n2096), .Y(n2570) );
  OR2X1_RVT U2555 ( .A1(n2007), .A2(n2572), .Y(n2096) );
  OR2X1_RVT U2556 ( .A1(n2007), .A2(n2187), .Y(n2565) );
  OR2X1_RVT U2557 ( .A1(n31), .A2(n12599), .Y(n2187) );
  OR2X1_RVT U2558 ( .A1(n2573), .A2(n1963), .Y(n2564) );
  AND4X1_RVT U2559 ( .A1(n2574), .A2(n2575), .A3(n2576), .A4(n2577), .Y(n2573)
         );
  OR2X1_RVT U2560 ( .A1(n12896), .A2(n2578), .Y(n2576) );
  OR2X1_RVT U2561 ( .A1(n2579), .A2(n12903), .Y(n2578) );
  AND2X1_RVT U2562 ( .A1(n2014), .A2(n2580), .Y(n2579) );
  OR2X1_RVT U2563 ( .A1(n12592), .A2(n2581), .Y(n2575) );
  OR2X1_RVT U2564 ( .A1(n2320), .A2(n1957), .Y(n2581) );
  OR2X1_RVT U2565 ( .A1(n1940), .A2(n1966), .Y(n2574) );
  OR2X1_RVT U2566 ( .A1(n12900), .A2(n2066), .Y(n1966) );
  OR2X1_RVT U2567 ( .A1(n2440), .A2(n2354), .Y(n2563) );
  OR2X1_RVT U2568 ( .A1(n12608), .A2(n1977), .Y(n2354) );
  AND4X1_RVT U2569 ( .A1(n2583), .A2(n2584), .A3(n2585), .A4(n2586), .Y(n2582)
         );
  AND4X1_RVT U2570 ( .A1(n2587), .A2(n2588), .A3(n2589), .A4(n2590), .Y(n2586)
         );
  AND4X1_RVT U2571 ( .A1(n2591), .A2(n2592), .A3(n2593), .A4(n2594), .Y(n2590)
         );
  OR2X1_RVT U2572 ( .A1(n2428), .A2(n2572), .Y(n2594) );
  OR2X1_RVT U2573 ( .A1(n12899), .A2(n12602), .Y(n2572) );
  OR2X1_RVT U2574 ( .A1(n12576), .A2(n12586), .Y(n2428) );
  OR2X1_RVT U2575 ( .A1(n2595), .A2(n2014), .Y(n2593) );
  AND2X1_RVT U2576 ( .A1(n1960), .A2(n2527), .Y(n2595) );
  OR2X1_RVT U2577 ( .A1(n31), .A2(n2596), .Y(n1960) );
  OR2X1_RVT U2578 ( .A1(n12576), .A2(n12896), .Y(n2596) );
  OR2X1_RVT U2579 ( .A1(n2597), .A2(n1942), .Y(n2592) );
  OR2X1_RVT U2580 ( .A1(n12590), .A2(n2103), .Y(n1942) );
  AND2X1_RVT U2581 ( .A1(n2078), .A2(n2598), .Y(n2597) );
  OR2X1_RVT U2582 ( .A1(n1957), .A2(n2159), .Y(n2598) );
  OR2X1_RVT U2583 ( .A1(n12594), .A2(n12582), .Y(n1957) );
  OR2X1_RVT U2584 ( .A1(n2203), .A2(n2599), .Y(n2078) );
  OR2X1_RVT U2585 ( .A1(n12907), .A2(n12597), .Y(n2599) );
  OR2X1_RVT U2586 ( .A1(n2600), .A2(n2001), .Y(n2591) );
  AND2X1_RVT U2587 ( .A1(n2398), .A2(n2601), .Y(n2600) );
  OR2X1_RVT U2588 ( .A1(n2602), .A2(n12896), .Y(n2601) );
  AND2X1_RVT U2589 ( .A1(n2057), .A2(n2410), .Y(n2602) );
  OR2X1_RVT U2590 ( .A1(n12904), .A2(n2019), .Y(n2410) );
  OR2X1_RVT U2591 ( .A1(n12603), .A2(n2603), .Y(n2398) );
  OR2X1_RVT U2592 ( .A1(n12909), .A2(n12905), .Y(n2603) );
  OR2X1_RVT U2593 ( .A1(n2604), .A2(n12581), .Y(n2589) );
  AND2X1_RVT U2594 ( .A1(n2605), .A2(n2606), .Y(n2604) );
  OR2X1_RVT U2595 ( .A1(n2607), .A2(n2103), .Y(n2606) );
  AND2X1_RVT U2596 ( .A1(n2168), .A2(n2608), .Y(n2607) );
  OR2X1_RVT U2597 ( .A1(n1959), .A2(n2081), .Y(n2605) );
  OR2X1_RVT U2598 ( .A1(n12595), .A2(n2017), .Y(n2081) );
  OR2X1_RVT U2599 ( .A1(n2609), .A2(n12905), .Y(n2588) );
  AND2X1_RVT U2600 ( .A1(n2173), .A2(n2332), .Y(n2609) );
  OR2X1_RVT U2601 ( .A1(n12593), .A2(n2610), .Y(n2332) );
  OR2X1_RVT U2602 ( .A1(n2013), .A2(n12582), .Y(n2610) );
  OR2X1_RVT U2603 ( .A1(n1959), .A2(n2440), .Y(n2173) );
  OR2X1_RVT U2604 ( .A1(n12582), .A2(n12597), .Y(n2440) );
  OR2X1_RVT U2605 ( .A1(n2611), .A2(n12579), .Y(n2587) );
  AND2X1_RVT U2606 ( .A1(n2213), .A2(n2612), .Y(n2611) );
  OR2X1_RVT U2607 ( .A1(n2427), .A2(n2007), .Y(n2612) );
  OR2X1_RVT U2608 ( .A1(n2066), .A2(n2548), .Y(n2213) );
  OR2X1_RVT U2609 ( .A1(n12904), .A2(n31), .Y(n2548) );
  AND2X1_RVT U2610 ( .A1(n12583), .A2(n12907), .Y(n2309) );
  AND4X1_RVT U2611 ( .A1(n2613), .A2(n2614), .A3(n2615), .A4(n2616), .Y(n2585)
         );
  AND4X1_RVT U2612 ( .A1(n2617), .A2(n2618), .A3(n2619), .A4(n2620), .Y(n2616)
         );
  OR2X1_RVT U2613 ( .A1(n2621), .A2(n12588), .Y(n2620) );
  AND2X1_RVT U2614 ( .A1(n2200), .A2(n2271), .Y(n2621) );
  OR2X1_RVT U2615 ( .A1(n2016), .A2(n2527), .Y(n2271) );
  OR2X1_RVT U2616 ( .A1(n12907), .A2(n2013), .Y(n2527) );
  OR2X1_RVT U2617 ( .A1(n12894), .A2(n12578), .Y(n2016) );
  OR2X1_RVT U2618 ( .A1(n12579), .A2(n2303), .Y(n2200) );
  OR2X1_RVT U2619 ( .A1(n12583), .A2(n12597), .Y(n2303) );
  OR2X1_RVT U2620 ( .A1(n2622), .A2(n12903), .Y(n2619) );
  AND2X1_RVT U2621 ( .A1(n2362), .A2(n2623), .Y(n2622) );
  OR2X1_RVT U2622 ( .A1(n2320), .A2(n2030), .Y(n2623) );
  OR2X1_RVT U2623 ( .A1(n2203), .A2(n2624), .Y(n2030) );
  OR2X1_RVT U2624 ( .A1(n12608), .A2(n12584), .Y(n2624) );
  OR2X1_RVT U2625 ( .A1(n12592), .A2(n2625), .Y(n2362) );
  OR2X1_RVT U2626 ( .A1(n2203), .A2(n1999), .Y(n2625) );
  OR2X1_RVT U2627 ( .A1(n2626), .A2(n12909), .Y(n2618) );
  AND2X1_RVT U2628 ( .A1(n2308), .A2(n2237), .Y(n2626) );
  OR2X1_RVT U2629 ( .A1(n2019), .A2(n2055), .Y(n2237) );
  OR2X1_RVT U2630 ( .A1(n12901), .A2(n2203), .Y(n2055) );
  OR2X1_RVT U2631 ( .A1(n2427), .A2(n2035), .Y(n2308) );
  OR2X1_RVT U2632 ( .A1(n12589), .A2(n12906), .Y(n2427) );
  OR2X1_RVT U2633 ( .A1(n2627), .A2(n2077), .Y(n2617) );
  AND2X1_RVT U2634 ( .A1(n2628), .A2(n2629), .Y(n2627) );
  OR2X1_RVT U2635 ( .A1(n1999), .A2(n2426), .Y(n2629) );
  OR2X1_RVT U2636 ( .A1(n12903), .A2(n39), .Y(n2426) );
  AND2X1_RVT U2637 ( .A1(n2630), .A2(n2294), .Y(n2628) );
  OR2X1_RVT U2638 ( .A1(n2007), .A2(n2631), .Y(n2294) );
  OR2X1_RVT U2639 ( .A1(n12605), .A2(n12584), .Y(n2631) );
  OR2X1_RVT U2640 ( .A1(n2063), .A2(n2000), .Y(n2615) );
  OR2X1_RVT U2641 ( .A1(n12896), .A2(n1959), .Y(n2063) );
  OR2X1_RVT U2642 ( .A1(n2632), .A2(n1963), .Y(n2614) );
  AND2X1_RVT U2643 ( .A1(n2633), .A2(n2144), .Y(n2632) );
  AND2X1_RVT U2644 ( .A1(n2634), .A2(n2635), .Y(n2144) );
  OR2X1_RVT U2645 ( .A1(n12593), .A2(n2168), .Y(n2635) );
  OR2X1_RVT U2646 ( .A1(n2066), .A2(n1940), .Y(n2634) );
  OR2X1_RVT U2647 ( .A1(n12578), .A2(n2013), .Y(n1940) );
  AND2X1_RVT U2648 ( .A1(n2636), .A2(n2330), .Y(n2633) );
  OR2X1_RVT U2649 ( .A1(n2097), .A2(n2580), .Y(n2330) );
  OR2X1_RVT U2650 ( .A1(n12898), .A2(n29), .Y(n2580) );
  OR2X1_RVT U2651 ( .A1(n1959), .A2(n2126), .Y(n2636) );
  OR2X1_RVT U2652 ( .A1(n12577), .A2(n2637), .Y(n2126) );
  OR2X1_RVT U2653 ( .A1(n12894), .A2(n12606), .Y(n2637) );
  OR2X1_RVT U2654 ( .A1(n2638), .A2(n12894), .Y(n2613) );
  AND4X1_RVT U2655 ( .A1(n2639), .A2(n2640), .A3(n2641), .A4(n2472), .Y(n2638)
         );
  OR2X1_RVT U2656 ( .A1(n2013), .A2(n2393), .Y(n2472) );
  OR2X1_RVT U2657 ( .A1(n12899), .A2(n12905), .Y(n2393) );
  OR2X1_RVT U2658 ( .A1(n2013), .A2(n2642), .Y(n2641) );
  OR2X1_RVT U2659 ( .A1(n12583), .A2(n12588), .Y(n2642) );
  OR2X1_RVT U2660 ( .A1(n12904), .A2(n1972), .Y(n2013) );
  OR2X1_RVT U2661 ( .A1(n2643), .A2(n2094), .Y(n2640) );
  OR2X1_RVT U2662 ( .A1(n12577), .A2(n1938), .Y(n2094) );
  AND2X1_RVT U2663 ( .A1(n2077), .A2(n2644), .Y(n2643) );
  OR2X1_RVT U2664 ( .A1(n12902), .A2(n1977), .Y(n2644) );
  OR2X1_RVT U2665 ( .A1(n12898), .A2(n12588), .Y(n2077) );
  OR2X1_RVT U2666 ( .A1(n12900), .A2(n2608), .Y(n2639) );
  OR2X1_RVT U2667 ( .A1(n12904), .A2(n2017), .Y(n2608) );
  OR2X1_RVT U2668 ( .A1(n1963), .A2(n29), .Y(n2017) );
  AND4X1_RVT U2669 ( .A1(n2645), .A2(n2646), .A3(n2647), .A4(n2648), .Y(n2584)
         );
  AND4X1_RVT U2670 ( .A1(n2649), .A2(n2650), .A3(n2651), .A4(n2652), .Y(n2648)
         );
  OR2X1_RVT U2671 ( .A1(n2035), .A2(n2162), .Y(n2652) );
  OR2X1_RVT U2672 ( .A1(n12590), .A2(n2057), .Y(n2162) );
  OR2X1_RVT U2673 ( .A1(n12594), .A2(n2203), .Y(n2035) );
  OR2X1_RVT U2674 ( .A1(n2022), .A2(n2498), .Y(n2651) );
  OR2X1_RVT U2675 ( .A1(n12908), .A2(n12577), .Y(n2498) );
  OR2X1_RVT U2676 ( .A1(n2088), .A2(n2014), .Y(n2022) );
  OR2X1_RVT U2677 ( .A1(n2007), .A2(n2034), .Y(n2650) );
  OR2X1_RVT U2678 ( .A1(n12586), .A2(n12599), .Y(n2034) );
  OR2X1_RVT U2679 ( .A1(n12576), .A2(n12895), .Y(n2007) );
  OR2X1_RVT U2680 ( .A1(n39), .A2(n2373), .Y(n2649) );
  OR2X1_RVT U2681 ( .A1(n12584), .A2(n2160), .Y(n2373) );
  OR2X1_RVT U2682 ( .A1(n1977), .A2(n2407), .Y(n2647) );
  OR2X1_RVT U2683 ( .A1(n39), .A2(n2653), .Y(n2407) );
  OR2X1_RVT U2684 ( .A1(n12901), .A2(n12597), .Y(n2653) );
  AND2X1_RVT U2685 ( .A1(n12578), .A2(n12581), .Y(n2437) );
  OR2X1_RVT U2686 ( .A1(n2019), .A2(n1967), .Y(n2646) );
  OR2X1_RVT U2687 ( .A1(n12606), .A2(n2654), .Y(n1967) );
  OR2X1_RVT U2688 ( .A1(n12902), .A2(n12894), .Y(n2654) );
  OR2X1_RVT U2689 ( .A1(n12583), .A2(n1999), .Y(n2019) );
  OR2X1_RVT U2690 ( .A1(n2066), .A2(n2630), .Y(n2645) );
  OR2X1_RVT U2691 ( .A1(n12579), .A2(n2021), .Y(n2630) );
  OR2X1_RVT U2692 ( .A1(n12904), .A2(n12905), .Y(n2021) );
  AND4X1_RVT U2693 ( .A1(n2655), .A2(n2132), .A3(n2656), .A4(n2657), .Y(n2583)
         );
  OR2X1_RVT U2694 ( .A1(n12583), .A2(n2577), .Y(n2657) );
  OR2X1_RVT U2695 ( .A1(n12900), .A2(n2127), .Y(n2577) );
  OR2X1_RVT U2696 ( .A1(n12581), .A2(n2168), .Y(n2127) );
  OR2X1_RVT U2697 ( .A1(n12576), .A2(n1994), .Y(n2168) );
  AND2X1_RVT U2698 ( .A1(n2658), .A2(n2659), .Y(n2656) );
  OR2X1_RVT U2699 ( .A1(n12605), .A2(n2497), .Y(n2659) );
  OR2X1_RVT U2700 ( .A1(n2066), .A2(n2159), .Y(n2497) );
  OR2X1_RVT U2701 ( .A1(n12583), .A2(n12577), .Y(n2159) );
  OR2X1_RVT U2702 ( .A1(n12578), .A2(n1955), .Y(n1994) );
  OR2X1_RVT U2703 ( .A1(n12907), .A2(n2228), .Y(n2658) );
  OR2X1_RVT U2704 ( .A1(n12602), .A2(n2262), .Y(n2228) );
  OR2X1_RVT U2705 ( .A1(n12899), .A2(n12894), .Y(n2262) );
  OR2X1_RVT U2706 ( .A1(n12897), .A2(n12594), .Y(n1938) );
  AND2X1_RVT U2707 ( .A1(n2660), .A2(n2661), .Y(n2132) );
  OR2X1_RVT U2708 ( .A1(n2014), .A2(n2000), .Y(n2661) );
  OR2X1_RVT U2709 ( .A1(n12906), .A2(n1972), .Y(n2000) );
  AND2X1_RVT U2710 ( .A1(n1999), .A2(n1963), .Y(n2052) );
  OR2X1_RVT U2711 ( .A1(n12589), .A2(n2066), .Y(n2014) );
  OR2X1_RVT U2712 ( .A1(n12895), .A2(n2103), .Y(n2066) );
  OR2X1_RVT U2713 ( .A1(n2662), .A2(n2057), .Y(n2660) );
  OR2X1_RVT U2714 ( .A1(n12583), .A2(n29), .Y(n2057) );
  AND2X1_RVT U2715 ( .A1(n12908), .A2(n12576), .Y(n2320) );
  OR2X1_RVT U2716 ( .A1(n12582), .A2(n2160), .Y(n2662) );
  OR2X1_RVT U2717 ( .A1(n12904), .A2(n12599), .Y(n2160) );
  AND2X1_RVT U2718 ( .A1(n2663), .A2(n2664), .Y(n2655) );
  OR2X1_RVT U2719 ( .A1(n1980), .A2(n2313), .Y(n2664) );
  OR2X1_RVT U2720 ( .A1(n12584), .A2(n2020), .Y(n2313) );
  OR2X1_RVT U2721 ( .A1(n12599), .A2(n2097), .Y(n2020) );
  OR2X1_RVT U2722 ( .A1(n12579), .A2(n12582), .Y(n2097) );
  OR2X1_RVT U2723 ( .A1(n12901), .A2(n12899), .Y(n1959) );
  OR2X1_RVT U2724 ( .A1(n12909), .A2(n12903), .Y(n1980) );
  XOR2X1_RVT U2725 ( .A1(key[116]), .A2(state[116]), .Y(n1955) );
  OR2X1_RVT U2726 ( .A1(n1972), .A2(n2101), .Y(n2663) );
  OR2X1_RVT U2727 ( .A1(n2203), .A2(n2394), .Y(n2101) );
  OR2X1_RVT U2728 ( .A1(n12586), .A2(n2001), .Y(n2394) );
  OR2X1_RVT U2729 ( .A1(n12902), .A2(n2103), .Y(n2001) );
  XOR2X1_RVT U2730 ( .A1(key[114]), .A2(state[114]), .Y(n2103) );
  XOR2X1_RVT U2731 ( .A1(key[115]), .A2(state[115]), .Y(n2037) );
  OR2X1_RVT U2732 ( .A1(n12907), .A2(n12584), .Y(n1977) );
  XOR2X1_RVT U2733 ( .A1(key[117]), .A2(state[117]), .Y(n1963) );
  XOR2X1_RVT U2734 ( .A1(key[118]), .A2(state[118]), .Y(n1999) );
  OR2X1_RVT U2735 ( .A1(n12897), .A2(n12582), .Y(n2203) );
  XOR2X1_RVT U2736 ( .A1(key[112]), .A2(state[112]), .Y(n1978) );
  XOR2X1_RVT U2737 ( .A1(key[113]), .A2(state[113]), .Y(n2088) );
  XOR2X1_RVT U2738 ( .A1(key[119]), .A2(state[119]), .Y(n1972) );
  AND4X1_RVT U2739 ( .A1(n2666), .A2(n2667), .A3(n2668), .A4(n2669), .Y(n2665)
         );
  AND4X1_RVT U2740 ( .A1(n2670), .A2(n2671), .A3(n2672), .A4(n2673), .Y(n2669)
         );
  AND4X1_RVT U2741 ( .A1(n2674), .A2(n2675), .A3(n2676), .A4(n2677), .Y(n2673)
         );
  OR2X1_RVT U2742 ( .A1(n12504), .A2(n2679), .Y(n2672) );
  OR2X1_RVT U2743 ( .A1(n2680), .A2(n2681), .Y(n2670) );
  OR2X1_RVT U2744 ( .A1(n12891), .A2(n2682), .Y(n2681) );
  AND4X1_RVT U2745 ( .A1(n2683), .A2(n2684), .A3(n2685), .A4(n2686), .Y(n2668)
         );
  OR2X1_RVT U2746 ( .A1(n2687), .A2(n12889), .Y(n2686) );
  AND2X1_RVT U2747 ( .A1(n2688), .A2(n2689), .Y(n2687) );
  AND2X1_RVT U2748 ( .A1(n2690), .A2(n2691), .Y(n2685) );
  OR2X1_RVT U2749 ( .A1(n2692), .A2(n51), .Y(n2691) );
  AND2X1_RVT U2750 ( .A1(n2693), .A2(n2694), .Y(n2692) );
  OR2X1_RVT U2751 ( .A1(n12495), .A2(n2696), .Y(n2694) );
  OR2X1_RVT U2752 ( .A1(n2682), .A2(n2697), .Y(n2693) );
  OR2X1_RVT U2753 ( .A1(n2698), .A2(n12501), .Y(n2690) );
  AND2X1_RVT U2754 ( .A1(n2700), .A2(n2701), .Y(n2698) );
  OR2X1_RVT U2755 ( .A1(n2702), .A2(n2703), .Y(n2684) );
  AND2X1_RVT U2756 ( .A1(n2704), .A2(n2705), .Y(n2702) );
  OR2X1_RVT U2757 ( .A1(n12496), .A2(n2706), .Y(n2705) );
  AND2X1_RVT U2758 ( .A1(n2707), .A2(n2708), .Y(n2704) );
  AND2X1_RVT U2759 ( .A1(n2709), .A2(n2710), .Y(n2683) );
  OR2X1_RVT U2760 ( .A1(n2711), .A2(n12478), .Y(n2710) );
  AND2X1_RVT U2761 ( .A1(n2713), .A2(n2714), .Y(n2711) );
  OR2X1_RVT U2762 ( .A1(n2715), .A2(n2716), .Y(n2714) );
  OR2X1_RVT U2763 ( .A1(n12487), .A2(n12482), .Y(n2716) );
  OR2X1_RVT U2764 ( .A1(n2719), .A2(n2720), .Y(n2709) );
  AND2X1_RVT U2765 ( .A1(n2721), .A2(n2722), .Y(n2719) );
  AND2X1_RVT U2766 ( .A1(n2723), .A2(n2724), .Y(n2721) );
  AND4X1_RVT U2767 ( .A1(n2725), .A2(n2726), .A3(n2727), .A4(n2728), .Y(n2667)
         );
  AND4X1_RVT U2768 ( .A1(n2729), .A2(n2730), .A3(n2731), .A4(n2732), .Y(n2728)
         );
  OR2X1_RVT U2769 ( .A1(n2733), .A2(n12507), .Y(n2732) );
  AND4X1_RVT U2770 ( .A1(n2735), .A2(n2736), .A3(n2737), .A4(n2738), .Y(n2733)
         );
  OR2X1_RVT U2771 ( .A1(n2739), .A2(n2706), .Y(n2738) );
  OR2X1_RVT U2772 ( .A1(n2740), .A2(n12493), .Y(n2737) );
  OR2X1_RVT U2773 ( .A1(n2742), .A2(n12484), .Y(n2731) );
  AND4X1_RVT U2774 ( .A1(n2743), .A2(n2744), .A3(n2745), .A4(n2746), .Y(n2742)
         );
  OR2X1_RVT U2775 ( .A1(n2747), .A2(n2748), .Y(n2746) );
  OR2X1_RVT U2776 ( .A1(n12501), .A2(n12496), .Y(n2748) );
  AND2X1_RVT U2777 ( .A1(n2749), .A2(n2750), .Y(n2745) );
  OR2X1_RVT U2778 ( .A1(n12893), .A2(n2751), .Y(n2744) );
  OR2X1_RVT U2779 ( .A1(n2752), .A2(n2753), .Y(n2743) );
  AND2X1_RVT U2780 ( .A1(n2754), .A2(n2755), .Y(n2752) );
  OR2X1_RVT U2781 ( .A1(n12501), .A2(n2756), .Y(n2755) );
  OR2X1_RVT U2782 ( .A1(n2689), .A2(n2757), .Y(n2730) );
  OR2X1_RVT U2783 ( .A1(n2756), .A2(n2758), .Y(n2729) );
  OR2X1_RVT U2784 ( .A1(n2759), .A2(n2760), .Y(n2727) );
  OR2X1_RVT U2785 ( .A1(n2761), .A2(n2754), .Y(n2726) );
  OR2X1_RVT U2786 ( .A1(n2762), .A2(n2763), .Y(n2725) );
  AND4X1_RVT U2787 ( .A1(n2764), .A2(n2765), .A3(n2766), .A4(n2767), .Y(n2666)
         );
  AND2X1_RVT U2788 ( .A1(n2768), .A2(n2769), .Y(n2767) );
  OR2X1_RVT U2789 ( .A1(n2753), .A2(n2770), .Y(n2769) );
  AND2X1_RVT U2790 ( .A1(n2771), .A2(n2772), .Y(n2768) );
  OR2X1_RVT U2791 ( .A1(n2773), .A2(n2696), .Y(n2772) );
  OR2X1_RVT U2792 ( .A1(n2697), .A2(n2774), .Y(n2771) );
  OR2X1_RVT U2793 ( .A1(n49), .A2(n2775), .Y(n2766) );
  OR2X1_RVT U2794 ( .A1(n2776), .A2(n12491), .Y(n2765) );
  OR2X1_RVT U2795 ( .A1(n12494), .A2(n2778), .Y(n2764) );
  AND4X1_RVT U2796 ( .A1(n2780), .A2(n2781), .A3(n2782), .A4(n2783), .Y(n2779)
         );
  AND4X1_RVT U2797 ( .A1(n2784), .A2(n2675), .A3(n2785), .A4(n2786), .Y(n2783)
         );
  AND4X1_RVT U2798 ( .A1(n2787), .A2(n2788), .A3(n2789), .A4(n2790), .Y(n2786)
         );
  OR2X1_RVT U2799 ( .A1(n2696), .A2(n2791), .Y(n2790) );
  OR2X1_RVT U2800 ( .A1(n2792), .A2(n12506), .Y(n2791) );
  OR2X1_RVT U2801 ( .A1(n2697), .A2(n2793), .Y(n2789) );
  OR2X1_RVT U2802 ( .A1(n49), .A2(n12490), .Y(n2793) );
  OR2X1_RVT U2803 ( .A1(n2794), .A2(n2740), .Y(n2788) );
  AND2X1_RVT U2804 ( .A1(n2751), .A2(n2795), .Y(n2794) );
  OR2X1_RVT U2805 ( .A1(n2796), .A2(n2797), .Y(n2787) );
  AND2X1_RVT U2806 ( .A1(n2798), .A2(n2799), .Y(n2796) );
  AND2X1_RVT U2807 ( .A1(n2800), .A2(n2801), .Y(n2785) );
  OR2X1_RVT U2808 ( .A1(n2747), .A2(n2802), .Y(n2801) );
  OR2X1_RVT U2809 ( .A1(n2803), .A2(n12891), .Y(n2802) );
  OR2X1_RVT U2810 ( .A1(n2804), .A2(n2805), .Y(n2800) );
  OR2X1_RVT U2811 ( .A1(n2806), .A2(n12495), .Y(n2805) );
  OR2X1_RVT U2812 ( .A1(n2682), .A2(n2807), .Y(n2675) );
  AND4X1_RVT U2813 ( .A1(n2808), .A2(n2809), .A3(n2810), .A4(n2811), .Y(n2782)
         );
  AND4X1_RVT U2814 ( .A1(n2812), .A2(n2813), .A3(n2814), .A4(n2815), .Y(n2811)
         );
  OR2X1_RVT U2815 ( .A1(n2816), .A2(n12509), .Y(n2815) );
  AND2X1_RVT U2816 ( .A1(n2818), .A2(n2819), .Y(n2816) );
  OR2X1_RVT U2817 ( .A1(n12478), .A2(n2697), .Y(n2819) );
  OR2X1_RVT U2818 ( .A1(n2820), .A2(n2699), .Y(n2814) );
  AND2X1_RVT U2819 ( .A1(n2821), .A2(n2822), .Y(n2820) );
  OR2X1_RVT U2820 ( .A1(n2823), .A2(n12890), .Y(n2813) );
  AND2X1_RVT U2821 ( .A1(n2824), .A2(n2825), .Y(n2823) );
  OR2X1_RVT U2822 ( .A1(n2826), .A2(n2775), .Y(n2825) );
  AND2X1_RVT U2823 ( .A1(n12509), .A2(n12493), .Y(n2826) );
  OR2X1_RVT U2824 ( .A1(n2827), .A2(n12479), .Y(n2812) );
  AND2X1_RVT U2825 ( .A1(n2829), .A2(n2830), .Y(n2827) );
  OR2X1_RVT U2826 ( .A1(n2831), .A2(n12485), .Y(n2810) );
  AND2X1_RVT U2827 ( .A1(n2832), .A2(n2833), .Y(n2831) );
  OR2X1_RVT U2828 ( .A1(n12493), .A2(n2834), .Y(n2833) );
  AND2X1_RVT U2829 ( .A1(n2835), .A2(n2836), .Y(n2832) );
  OR2X1_RVT U2830 ( .A1(n2837), .A2(n2838), .Y(n2835) );
  OR2X1_RVT U2831 ( .A1(n2682), .A2(n2753), .Y(n2838) );
  OR2X1_RVT U2832 ( .A1(n2839), .A2(n12887), .Y(n2809) );
  AND2X1_RVT U2833 ( .A1(n2840), .A2(n2841), .Y(n2839) );
  OR2X1_RVT U2834 ( .A1(n2842), .A2(n2843), .Y(n2808) );
  AND2X1_RVT U2835 ( .A1(n2844), .A2(n2845), .Y(n2842) );
  AND2X1_RVT U2836 ( .A1(n2846), .A2(n2847), .Y(n2844) );
  OR2X1_RVT U2837 ( .A1(n51), .A2(n2775), .Y(n2847) );
  OR2X1_RVT U2838 ( .A1(n12503), .A2(n2740), .Y(n2846) );
  AND4X1_RVT U2839 ( .A1(n2848), .A2(n2849), .A3(n2850), .A4(n2851), .Y(n2781)
         );
  AND4X1_RVT U2840 ( .A1(n2852), .A2(n2853), .A3(n2854), .A4(n2855), .Y(n2851)
         );
  OR2X1_RVT U2841 ( .A1(n2775), .A2(n2774), .Y(n2855) );
  OR2X1_RVT U2842 ( .A1(n2706), .A2(n2856), .Y(n2854) );
  OR2X1_RVT U2843 ( .A1(n2739), .A2(n2857), .Y(n2853) );
  OR2X1_RVT U2844 ( .A1(n2682), .A2(n2858), .Y(n2852) );
  AND2X1_RVT U2845 ( .A1(n2859), .A2(n2860), .Y(n2850) );
  OR2X1_RVT U2846 ( .A1(n12504), .A2(n2861), .Y(n2860) );
  OR2X1_RVT U2847 ( .A1(n12483), .A2(n2758), .Y(n2859) );
  OR2X1_RVT U2848 ( .A1(n2862), .A2(n2717), .Y(n2849) );
  AND4X1_RVT U2849 ( .A1(n2863), .A2(n2864), .A3(n2865), .A4(n2866), .Y(n2862)
         );
  OR2X1_RVT U2850 ( .A1(n2867), .A2(n2682), .Y(n2865) );
  OR2X1_RVT U2851 ( .A1(n12879), .A2(n2868), .Y(n2864) );
  OR2X1_RVT U2852 ( .A1(n2869), .A2(n12887), .Y(n2863) );
  AND2X1_RVT U2853 ( .A1(n2760), .A2(n2870), .Y(n2869) );
  OR2X1_RVT U2854 ( .A1(n2762), .A2(n2871), .Y(n2848) );
  AND4X1_RVT U2855 ( .A1(n2872), .A2(n2873), .A3(n2874), .A4(n2875), .Y(n2780)
         );
  AND4X1_RVT U2856 ( .A1(n2876), .A2(n2877), .A3(n2878), .A4(n2879), .Y(n2875)
         );
  OR2X1_RVT U2857 ( .A1(n12883), .A2(n2880), .Y(n2879) );
  OR2X1_RVT U2858 ( .A1(n12884), .A2(n2881), .Y(n2878) );
  OR2X1_RVT U2859 ( .A1(n12881), .A2(n2882), .Y(n2877) );
  OR2X1_RVT U2860 ( .A1(n12477), .A2(n2883), .Y(n2876) );
  OR2X1_RVT U2861 ( .A1(n2884), .A2(n12484), .Y(n2873) );
  AND4X1_RVT U2862 ( .A1(n2886), .A2(n2887), .A3(n2888), .A4(n2889), .Y(n2885)
         );
  AND4X1_RVT U2863 ( .A1(n2890), .A2(n2891), .A3(n2892), .A4(n2893), .Y(n2889)
         );
  AND4X1_RVT U2864 ( .A1(n2894), .A2(n2671), .A3(n2841), .A4(n2895), .Y(n2893)
         );
  OR2X1_RVT U2865 ( .A1(n2896), .A2(n12878), .Y(n2671) );
  AND2X1_RVT U2866 ( .A1(n2897), .A2(n2898), .Y(n2896) );
  OR2X1_RVT U2867 ( .A1(n2715), .A2(n2899), .Y(n2898) );
  OR2X1_RVT U2868 ( .A1(n2900), .A2(n2797), .Y(n2897) );
  OR2X1_RVT U2869 ( .A1(n2901), .A2(n2756), .Y(n2894) );
  AND2X1_RVT U2870 ( .A1(n2902), .A2(n2903), .Y(n2901) );
  OR2X1_RVT U2871 ( .A1(n12883), .A2(n2740), .Y(n2903) );
  OR2X1_RVT U2872 ( .A1(n2904), .A2(n2699), .Y(n2892) );
  AND2X1_RVT U2873 ( .A1(n2905), .A2(n2906), .Y(n2904) );
  OR2X1_RVT U2874 ( .A1(n2907), .A2(n12889), .Y(n2906) );
  AND2X1_RVT U2875 ( .A1(n2747), .A2(n2908), .Y(n2907) );
  OR2X1_RVT U2876 ( .A1(n2909), .A2(n12504), .Y(n2891) );
  AND2X1_RVT U2877 ( .A1(n2910), .A2(n2911), .Y(n2909) );
  OR2X1_RVT U2878 ( .A1(n2740), .A2(n2706), .Y(n2911) );
  OR2X1_RVT U2879 ( .A1(n2912), .A2(n12487), .Y(n2890) );
  AND2X1_RVT U2880 ( .A1(n2824), .A2(n2913), .Y(n2912) );
  OR2X1_RVT U2881 ( .A1(n2753), .A2(n2914), .Y(n2824) );
  AND4X1_RVT U2882 ( .A1(n2915), .A2(n2916), .A3(n2917), .A4(n2918), .Y(n2888)
         );
  OR2X1_RVT U2883 ( .A1(n2919), .A2(n12494), .Y(n2918) );
  AND2X1_RVT U2884 ( .A1(n2920), .A2(n2921), .Y(n2919) );
  OR2X1_RVT U2885 ( .A1(n2797), .A2(n2697), .Y(n2921) );
  AND2X1_RVT U2886 ( .A1(n2922), .A2(n2923), .Y(n2920) );
  OR2X1_RVT U2887 ( .A1(n2837), .A2(n2899), .Y(n2922) );
  AND2X1_RVT U2888 ( .A1(n2924), .A2(n2925), .Y(n2917) );
  OR2X1_RVT U2889 ( .A1(n2926), .A2(n2828), .Y(n2925) );
  AND2X1_RVT U2890 ( .A1(n2927), .A2(n2736), .Y(n2926) );
  OR2X1_RVT U2891 ( .A1(n2682), .A2(n2797), .Y(n2736) );
  OR2X1_RVT U2892 ( .A1(n2928), .A2(n51), .Y(n2924) );
  AND2X1_RVT U2893 ( .A1(n2929), .A2(n2930), .Y(n2928) );
  OR2X1_RVT U2894 ( .A1(n2931), .A2(n12496), .Y(n2930) );
  AND2X1_RVT U2895 ( .A1(n2932), .A2(n2933), .Y(n2931) );
  OR2X1_RVT U2896 ( .A1(n12491), .A2(n2747), .Y(n2933) );
  OR2X1_RVT U2897 ( .A1(n12893), .A2(n12493), .Y(n2932) );
  AND2X1_RVT U2898 ( .A1(n2798), .A2(n2908), .Y(n2929) );
  OR2X1_RVT U2899 ( .A1(n2828), .A2(n2934), .Y(n2798) );
  OR2X1_RVT U2900 ( .A1(n12888), .A2(n12884), .Y(n2934) );
  OR2X1_RVT U2901 ( .A1(n2935), .A2(n2817), .Y(n2916) );
  AND4X1_RVT U2902 ( .A1(n2776), .A2(n2936), .A3(n2937), .A4(n2938), .Y(n2935)
         );
  OR2X1_RVT U2903 ( .A1(n12495), .A2(n2797), .Y(n2938) );
  AND2X1_RVT U2904 ( .A1(n2939), .A2(n2940), .Y(n2937) );
  OR2X1_RVT U2905 ( .A1(n12893), .A2(n12504), .Y(n2936) );
  AND2X1_RVT U2906 ( .A1(n2941), .A2(n2942), .Y(n2776) );
  OR2X1_RVT U2907 ( .A1(n2943), .A2(n49), .Y(n2942) );
  OR2X1_RVT U2908 ( .A1(n2740), .A2(n12878), .Y(n2941) );
  AND2X1_RVT U2909 ( .A1(n2944), .A2(n2945), .Y(n2915) );
  OR2X1_RVT U2910 ( .A1(n2946), .A2(n12880), .Y(n2945) );
  AND2X1_RVT U2911 ( .A1(n2947), .A2(n2948), .Y(n2946) );
  OR2X1_RVT U2912 ( .A1(n2949), .A2(n12498), .Y(n2948) );
  AND2X1_RVT U2913 ( .A1(n2950), .A2(n2951), .Y(n2949) );
  AND2X1_RVT U2914 ( .A1(n2952), .A2(n2953), .Y(n2947) );
  OR2X1_RVT U2915 ( .A1(n2954), .A2(n12507), .Y(n2944) );
  AND4X1_RVT U2916 ( .A1(n2955), .A2(n2956), .A3(n2957), .A4(n2958), .Y(n2954)
         );
  OR2X1_RVT U2917 ( .A1(n12892), .A2(n2959), .Y(n2957) );
  OR2X1_RVT U2918 ( .A1(n49), .A2(n2754), .Y(n2956) );
  OR2X1_RVT U2919 ( .A1(n2843), .A2(n2797), .Y(n2955) );
  AND4X1_RVT U2920 ( .A1(n2960), .A2(n2961), .A3(n2962), .A4(n2963), .Y(n2887)
         );
  AND2X1_RVT U2921 ( .A1(n2964), .A2(n2807), .Y(n2963) );
  OR2X1_RVT U2922 ( .A1(n12482), .A2(n2773), .Y(n2807) );
  AND2X1_RVT U2923 ( .A1(n2965), .A2(n2966), .Y(n2964) );
  OR2X1_RVT U2924 ( .A1(n2967), .A2(n2722), .Y(n2966) );
  OR2X1_RVT U2925 ( .A1(n2774), .A2(n2834), .Y(n2965) );
  OR2X1_RVT U2926 ( .A1(n49), .A2(n2968), .Y(n2962) );
  OR2X1_RVT U2927 ( .A1(n12891), .A2(n2969), .Y(n2961) );
  OR2X1_RVT U2928 ( .A1(n2843), .A2(n2970), .Y(n2960) );
  AND4X1_RVT U2929 ( .A1(n2971), .A2(n2972), .A3(n2973), .A4(n2974), .Y(n2886)
         );
  AND2X1_RVT U2930 ( .A1(n2975), .A2(n2976), .Y(n2974) );
  OR2X1_RVT U2931 ( .A1(n12477), .A2(n2977), .Y(n2976) );
  AND2X1_RVT U2932 ( .A1(n2978), .A2(n2979), .Y(n2975) );
  OR2X1_RVT U2933 ( .A1(n2739), .A2(n2749), .Y(n2979) );
  OR2X1_RVT U2934 ( .A1(n12498), .A2(n2799), .Y(n2749) );
  OR2X1_RVT U2935 ( .A1(n12484), .A2(n2980), .Y(n2978) );
  OR2X1_RVT U2936 ( .A1(n2720), .A2(n2713), .Y(n2973) );
  OR2X1_RVT U2937 ( .A1(n2806), .A2(n2981), .Y(n2713) );
  OR2X1_RVT U2938 ( .A1(n12887), .A2(n2982), .Y(n2972) );
  OR2X1_RVT U2939 ( .A1(n12496), .A2(n2840), .Y(n2971) );
  OR2X1_RVT U2940 ( .A1(n12878), .A2(n2902), .Y(n2840) );
  AND4X1_RVT U2941 ( .A1(n2984), .A2(n2985), .A3(n2986), .A4(n2987), .Y(n2983)
         );
  AND4X1_RVT U2942 ( .A1(n2988), .A2(n2989), .A3(n2990), .A4(n2991), .Y(n2987)
         );
  OR2X1_RVT U2943 ( .A1(n59), .A2(n2992), .Y(n2991) );
  OR2X1_RVT U2944 ( .A1(n2993), .A2(n12509), .Y(n2992) );
  AND2X1_RVT U2945 ( .A1(n12498), .A2(n2759), .Y(n2993) );
  AND2X1_RVT U2946 ( .A1(n2674), .A2(n2994), .Y(n2990) );
  OR2X1_RVT U2947 ( .A1(n12487), .A2(n2995), .Y(n2674) );
  OR2X1_RVT U2948 ( .A1(n59), .A2(n2753), .Y(n2995) );
  OR2X1_RVT U2949 ( .A1(n2996), .A2(n2682), .Y(n2989) );
  AND2X1_RVT U2950 ( .A1(n2997), .A2(n2998), .Y(n2996) );
  AND2X1_RVT U2951 ( .A1(n2999), .A2(n3000), .Y(n2988) );
  OR2X1_RVT U2952 ( .A1(n3001), .A2(n3002), .Y(n3000) );
  AND2X1_RVT U2953 ( .A1(n3003), .A2(n2763), .Y(n3001) );
  OR2X1_RVT U2954 ( .A1(n3004), .A2(n2754), .Y(n2999) );
  AND2X1_RVT U2955 ( .A1(n2939), .A2(n2773), .Y(n3004) );
  OR2X1_RVT U2956 ( .A1(n12485), .A2(n3005), .Y(n2939) );
  OR2X1_RVT U2957 ( .A1(n12893), .A2(n12495), .Y(n3005) );
  AND4X1_RVT U2958 ( .A1(n3006), .A2(n3007), .A3(n3008), .A4(n3009), .Y(n2986)
         );
  OR2X1_RVT U2959 ( .A1(n3010), .A2(n12883), .Y(n3009) );
  AND2X1_RVT U2960 ( .A1(n2822), .A2(n3011), .Y(n3010) );
  OR2X1_RVT U2961 ( .A1(n12891), .A2(n2867), .Y(n2822) );
  AND2X1_RVT U2962 ( .A1(n3012), .A2(n3013), .Y(n3008) );
  OR2X1_RVT U2963 ( .A1(n3014), .A2(n12881), .Y(n3013) );
  AND2X1_RVT U2964 ( .A1(n3015), .A2(n3016), .Y(n3014) );
  OR2X1_RVT U2965 ( .A1(n2717), .A2(n2959), .Y(n3016) );
  OR2X1_RVT U2966 ( .A1(n3017), .A2(n12879), .Y(n3012) );
  AND2X1_RVT U2967 ( .A1(n3018), .A2(n3019), .Y(n3017) );
  OR2X1_RVT U2968 ( .A1(n3020), .A2(n12498), .Y(n3007) );
  AND2X1_RVT U2969 ( .A1(n3021), .A2(n3022), .Y(n3020) );
  AND2X1_RVT U2970 ( .A1(n3023), .A2(n3024), .Y(n3021) );
  AND2X1_RVT U2971 ( .A1(n3025), .A2(n3026), .Y(n3006) );
  OR2X1_RVT U2972 ( .A1(n3027), .A2(n2943), .Y(n3026) );
  AND2X1_RVT U2973 ( .A1(n3028), .A2(n2774), .Y(n3027) );
  AND2X1_RVT U2974 ( .A1(n3029), .A2(n3030), .Y(n3028) );
  OR2X1_RVT U2975 ( .A1(n3031), .A2(n12501), .Y(n3025) );
  AND2X1_RVT U2976 ( .A1(n3032), .A2(n3033), .Y(n3031) );
  OR2X1_RVT U2977 ( .A1(n12890), .A2(n12503), .Y(n3033) );
  AND2X1_RVT U2978 ( .A1(n2763), .A2(n3034), .Y(n3032) );
  AND4X1_RVT U2979 ( .A1(n3035), .A2(n3036), .A3(n3037), .A4(n3038), .Y(n2985)
         );
  AND2X1_RVT U2980 ( .A1(n3039), .A2(n3040), .Y(n3038) );
  OR2X1_RVT U2981 ( .A1(n2756), .A2(n2830), .Y(n3040) );
  OR2X1_RVT U2982 ( .A1(n12885), .A2(n2763), .Y(n2830) );
  AND2X1_RVT U2983 ( .A1(n3041), .A2(n3042), .Y(n3039) );
  OR2X1_RVT U2984 ( .A1(n2908), .A2(n2722), .Y(n3042) );
  OR2X1_RVT U2985 ( .A1(n12892), .A2(n12494), .Y(n2722) );
  OR2X1_RVT U2986 ( .A1(n2806), .A2(n2856), .Y(n3041) );
  OR2X1_RVT U2987 ( .A1(n12880), .A2(n3043), .Y(n2856) );
  OR2X1_RVT U2988 ( .A1(n3044), .A2(n12477), .Y(n3037) );
  AND4X1_RVT U2989 ( .A1(n3045), .A2(n3046), .A3(n3047), .A4(n3048), .Y(n3044)
         );
  OR2X1_RVT U2990 ( .A1(n2981), .A2(n2754), .Y(n3047) );
  OR2X1_RVT U2991 ( .A1(n3049), .A2(n2751), .Y(n3046) );
  OR2X1_RVT U2992 ( .A1(n12889), .A2(n2706), .Y(n3045) );
  OR2X1_RVT U2993 ( .A1(n3050), .A2(n12478), .Y(n3036) );
  AND2X1_RVT U2994 ( .A1(n3051), .A2(n3052), .Y(n3050) );
  OR2X1_RVT U2995 ( .A1(n2981), .A2(n2706), .Y(n3052) );
  AND2X1_RVT U2996 ( .A1(n3053), .A2(n2982), .Y(n3051) );
  OR2X1_RVT U2997 ( .A1(n2754), .A2(n3054), .Y(n2982) );
  OR2X1_RVT U2998 ( .A1(n12880), .A2(n12892), .Y(n3054) );
  OR2X1_RVT U2999 ( .A1(n3055), .A2(n12485), .Y(n3035) );
  AND4X1_RVT U3000 ( .A1(n3056), .A2(n2969), .A3(n2778), .A4(n2750), .Y(n3055)
         );
  OR2X1_RVT U3001 ( .A1(n2775), .A2(n3057), .Y(n2750) );
  OR2X1_RVT U3002 ( .A1(n12882), .A2(n2712), .Y(n3057) );
  OR2X1_RVT U3003 ( .A1(n2837), .A2(n2871), .Y(n2778) );
  OR2X1_RVT U3004 ( .A1(n2756), .A2(n3058), .Y(n2969) );
  OR2X1_RVT U3005 ( .A1(n12509), .A2(n12478), .Y(n3058) );
  OR2X1_RVT U3006 ( .A1(n2715), .A2(n3059), .Y(n3056) );
  OR2X1_RVT U3007 ( .A1(n3060), .A2(n12483), .Y(n3059) );
  AND4X1_RVT U3008 ( .A1(n3061), .A2(n3062), .A3(n3063), .A4(n3064), .Y(n2984)
         );
  AND2X1_RVT U3009 ( .A1(n3065), .A2(n3066), .Y(n3064) );
  AND2X1_RVT U3010 ( .A1(n3067), .A2(n3068), .Y(n3065) );
  OR2X1_RVT U3011 ( .A1(n2747), .A2(n3022), .Y(n3068) );
  OR2X1_RVT U3012 ( .A1(n2759), .A2(n3069), .Y(n3022) );
  OR2X1_RVT U3013 ( .A1(n12881), .A2(n12883), .Y(n3069) );
  OR2X1_RVT U3014 ( .A1(n12888), .A2(n3070), .Y(n3067) );
  OR2X1_RVT U3015 ( .A1(n12494), .A2(n3071), .Y(n3063) );
  OR2X1_RVT U3016 ( .A1(n12891), .A2(n3072), .Y(n3062) );
  OR2X1_RVT U3017 ( .A1(n2759), .A2(n3073), .Y(n3061) );
  AND4X1_RVT U3018 ( .A1(n3075), .A2(n3076), .A3(n3077), .A4(n3078), .Y(n3074)
         );
  AND4X1_RVT U3019 ( .A1(n3079), .A2(n3080), .A3(n3081), .A4(n3082), .Y(n3078)
         );
  AND4X1_RVT U3020 ( .A1(n3083), .A2(n3084), .A3(n2676), .A4(n3085), .Y(n3082)
         );
  OR2X1_RVT U3021 ( .A1(n2817), .A2(n3086), .Y(n2676) );
  OR2X1_RVT U3022 ( .A1(n2908), .A2(n51), .Y(n3086) );
  OR2X1_RVT U3023 ( .A1(n2680), .A2(n3087), .Y(n3084) );
  OR2X1_RVT U3024 ( .A1(n12886), .A2(n12889), .Y(n3087) );
  OR2X1_RVT U3025 ( .A1(n2943), .A2(n3088), .Y(n3083) );
  OR2X1_RVT U3026 ( .A1(n3089), .A2(n2717), .Y(n3088) );
  AND2X1_RVT U3027 ( .A1(n12498), .A2(n2817), .Y(n3089) );
  OR2X1_RVT U3028 ( .A1(n3090), .A2(n12504), .Y(n3081) );
  AND2X1_RVT U3029 ( .A1(n2958), .A2(n3030), .Y(n3090) );
  OR2X1_RVT U3030 ( .A1(n51), .A2(n3091), .Y(n3030) );
  OR2X1_RVT U3031 ( .A1(n12477), .A2(n12885), .Y(n3091) );
  OR2X1_RVT U3032 ( .A1(n2747), .A2(n3092), .Y(n2958) );
  OR2X1_RVT U3033 ( .A1(n12883), .A2(n2739), .Y(n3092) );
  OR2X1_RVT U3034 ( .A1(n3093), .A2(n2697), .Y(n3080) );
  AND2X1_RVT U3035 ( .A1(n3094), .A2(n2902), .Y(n3093) );
  OR2X1_RVT U3036 ( .A1(n2803), .A2(n2797), .Y(n3079) );
  AND4X1_RVT U3037 ( .A1(n3095), .A2(n3096), .A3(n3097), .A4(n3098), .Y(n3077)
         );
  AND2X1_RVT U3038 ( .A1(n3099), .A2(n3100), .Y(n3098) );
  OR2X1_RVT U3039 ( .A1(n3101), .A2(n12498), .Y(n3100) );
  AND2X1_RVT U3040 ( .A1(n3102), .A2(n2770), .Y(n3101) );
  AND2X1_RVT U3041 ( .A1(n3103), .A2(n3104), .Y(n3099) );
  OR2X1_RVT U3042 ( .A1(n3105), .A2(n2753), .Y(n3104) );
  AND2X1_RVT U3043 ( .A1(n2724), .A2(n2696), .Y(n3105) );
  OR2X1_RVT U3044 ( .A1(n12891), .A2(n2795), .Y(n2724) );
  OR2X1_RVT U3045 ( .A1(n3106), .A2(n2806), .Y(n3103) );
  AND2X1_RVT U3046 ( .A1(n2998), .A2(n3107), .Y(n3106) );
  OR2X1_RVT U3047 ( .A1(n12892), .A2(n2834), .Y(n2998) );
  OR2X1_RVT U3048 ( .A1(n3108), .A2(n12883), .Y(n3097) );
  AND2X1_RVT U3049 ( .A1(n2701), .A2(n3109), .Y(n3108) );
  OR2X1_RVT U3050 ( .A1(n2837), .A2(n2761), .Y(n3109) );
  OR2X1_RVT U3051 ( .A1(n2740), .A2(n2943), .Y(n2701) );
  OR2X1_RVT U3052 ( .A1(n3110), .A2(n49), .Y(n3096) );
  AND2X1_RVT U3053 ( .A1(n2751), .A2(n3111), .Y(n3110) );
  OR2X1_RVT U3054 ( .A1(n3112), .A2(n12482), .Y(n3111) );
  AND2X1_RVT U3055 ( .A1(n3113), .A2(n3114), .Y(n3112) );
  OR2X1_RVT U3056 ( .A1(n12884), .A2(n2734), .Y(n3114) );
  OR2X1_RVT U3057 ( .A1(n12509), .A2(n2837), .Y(n2751) );
  OR2X1_RVT U3058 ( .A1(n3115), .A2(n2821), .Y(n3095) );
  AND2X1_RVT U3059 ( .A1(n2754), .A2(n2799), .Y(n3115) );
  OR2X1_RVT U3060 ( .A1(n12880), .A2(n2682), .Y(n2799) );
  AND4X1_RVT U3061 ( .A1(n3116), .A2(n3117), .A3(n3118), .A4(n3119), .Y(n3076)
         );
  AND4X1_RVT U3062 ( .A1(n3120), .A2(n3121), .A3(n3122), .A4(n3123), .Y(n3119)
         );
  OR2X1_RVT U3063 ( .A1(n3124), .A2(n12891), .Y(n3123) );
  AND2X1_RVT U3064 ( .A1(n2857), .A2(n3125), .Y(n3124) );
  OR2X1_RVT U3065 ( .A1(n12506), .A2(n2706), .Y(n3125) );
  OR2X1_RVT U3066 ( .A1(n3126), .A2(n2699), .Y(n3122) );
  AND2X1_RVT U3067 ( .A1(n3127), .A2(n3128), .Y(n3126) );
  OR2X1_RVT U3068 ( .A1(n3129), .A2(n2734), .Y(n3128) );
  AND2X1_RVT U3069 ( .A1(n2759), .A2(n2747), .Y(n3129) );
  AND2X1_RVT U3070 ( .A1(n2761), .A2(n3003), .Y(n3127) );
  OR2X1_RVT U3071 ( .A1(n12507), .A2(n2899), .Y(n3003) );
  OR2X1_RVT U3072 ( .A1(n3130), .A2(n12496), .Y(n3121) );
  AND2X1_RVT U3073 ( .A1(n3131), .A2(n3132), .Y(n3130) );
  OR2X1_RVT U3074 ( .A1(n2747), .A2(n3133), .Y(n3132) );
  AND2X1_RVT U3075 ( .A1(n2829), .A2(n3023), .Y(n3131) );
  OR2X1_RVT U3076 ( .A1(n2739), .A2(n2914), .Y(n3023) );
  OR2X1_RVT U3077 ( .A1(n2712), .A2(n3134), .Y(n2829) );
  OR2X1_RVT U3078 ( .A1(n3135), .A2(n2682), .Y(n3120) );
  AND4X1_RVT U3079 ( .A1(n3136), .A2(n3137), .A3(n3138), .A4(n3071), .Y(n3135)
         );
  OR2X1_RVT U3080 ( .A1(n2775), .A2(n3139), .Y(n3071) );
  OR2X1_RVT U3081 ( .A1(n12477), .A2(n2739), .Y(n3139) );
  OR2X1_RVT U3082 ( .A1(n12888), .A2(n2981), .Y(n3137) );
  OR2X1_RVT U3083 ( .A1(n2740), .A2(n2837), .Y(n3136) );
  OR2X1_RVT U3084 ( .A1(n2908), .A2(n2950), .Y(n3118) );
  OR2X1_RVT U3085 ( .A1(n3140), .A2(n12480), .Y(n3117) );
  AND4X1_RVT U3086 ( .A1(n3141), .A2(n3142), .A3(n2784), .A4(n2882), .Y(n3140)
         );
  OR2X1_RVT U3087 ( .A1(n2706), .A2(n2871), .Y(n2882) );
  OR2X1_RVT U3088 ( .A1(n12888), .A2(n49), .Y(n2871) );
  OR2X1_RVT U3089 ( .A1(n2699), .A2(n2763), .Y(n2784) );
  OR2X1_RVT U3090 ( .A1(n12880), .A2(n3134), .Y(n3116) );
  AND4X1_RVT U3091 ( .A1(n3143), .A2(n3144), .A3(n3145), .A4(n3146), .Y(n3075)
         );
  OR2X1_RVT U3092 ( .A1(n12485), .A2(n3147), .Y(n3146) );
  AND2X1_RVT U3093 ( .A1(n3148), .A2(n3149), .Y(n3145) );
  OR2X1_RVT U3094 ( .A1(n12506), .A2(n2902), .Y(n3149) );
  OR2X1_RVT U3095 ( .A1(n2689), .A2(n2763), .Y(n3148) );
  OR2X1_RVT U3096 ( .A1(n51), .A2(n2720), .Y(n2763) );
  OR2X1_RVT U3097 ( .A1(n12509), .A2(n2881), .Y(n3144) );
  OR2X1_RVT U3098 ( .A1(n2756), .A2(n3150), .Y(n2881) );
  AND2X1_RVT U3099 ( .A1(n3151), .A2(n3152), .Y(n3143) );
  OR2X1_RVT U3100 ( .A1(n12478), .A2(n3153), .Y(n3152) );
  OR2X1_RVT U3101 ( .A1(n2759), .A2(n2708), .Y(n3151) );
  OR2X1_RVT U3102 ( .A1(n2682), .A2(n2967), .Y(n2708) );
  AND4X1_RVT U3103 ( .A1(n3155), .A2(n3156), .A3(n3157), .A4(n3158), .Y(n3154)
         );
  AND4X1_RVT U3104 ( .A1(n3159), .A2(n3160), .A3(n3161), .A4(n3162), .Y(n3158)
         );
  AND4X1_RVT U3105 ( .A1(n2895), .A2(n3085), .A3(n3163), .A4(n3164), .Y(n3162)
         );
  OR2X1_RVT U3106 ( .A1(n3165), .A2(n3166), .Y(n3085) );
  OR2X1_RVT U3107 ( .A1(n2680), .A2(n2950), .Y(n2895) );
  OR2X1_RVT U3108 ( .A1(n12889), .A2(n12494), .Y(n2950) );
  AND4X1_RVT U3109 ( .A1(n3153), .A2(n3019), .A3(n3142), .A4(n2677), .Y(n3161)
         );
  OR2X1_RVT U3110 ( .A1(n3167), .A2(n2867), .Y(n2677) );
  OR2X1_RVT U3111 ( .A1(n2682), .A2(n3168), .Y(n3142) );
  OR2X1_RVT U3112 ( .A1(n2715), .A2(n49), .Y(n3019) );
  OR2X1_RVT U3113 ( .A1(n2706), .A2(n3169), .Y(n3153) );
  OR2X1_RVT U3114 ( .A1(n12484), .A2(n12504), .Y(n3169) );
  AND4X1_RVT U3115 ( .A1(n3170), .A2(n3171), .A3(n3172), .A4(n3173), .Y(n3160)
         );
  OR2X1_RVT U3116 ( .A1(n2959), .A2(n3174), .Y(n3173) );
  OR2X1_RVT U3117 ( .A1(n12504), .A2(n2739), .Y(n3174) );
  OR2X1_RVT U3118 ( .A1(n2868), .A2(n3175), .Y(n3172) );
  OR2X1_RVT U3119 ( .A1(n12890), .A2(n2756), .Y(n3175) );
  OR2X1_RVT U3120 ( .A1(n3094), .A2(n3176), .Y(n3171) );
  OR2X1_RVT U3121 ( .A1(n3177), .A2(n2753), .Y(n3176) );
  OR2X1_RVT U3122 ( .A1(n12501), .A2(n3178), .Y(n3170) );
  OR2X1_RVT U3123 ( .A1(n3179), .A2(n12484), .Y(n3178) );
  AND2X1_RVT U3124 ( .A1(n2967), .A2(n3180), .Y(n3179) );
  AND2X1_RVT U3125 ( .A1(n3181), .A2(n3182), .Y(n3159) );
  OR2X1_RVT U3126 ( .A1(n3183), .A2(n2734), .Y(n3182) );
  AND2X1_RVT U3127 ( .A1(n3184), .A2(n3185), .Y(n3183) );
  OR2X1_RVT U3128 ( .A1(n12483), .A2(n2927), .Y(n3185) );
  OR2X1_RVT U3129 ( .A1(n12487), .A2(n3002), .Y(n3184) );
  AND2X1_RVT U3130 ( .A1(n3186), .A2(n3187), .Y(n3181) );
  OR2X1_RVT U3131 ( .A1(n3188), .A2(n2773), .Y(n3187) );
  AND2X1_RVT U3132 ( .A1(n3189), .A2(n3190), .Y(n3188) );
  OR2X1_RVT U3133 ( .A1(n12490), .A2(n59), .Y(n3190) );
  NAND2X1_RVT U3134 ( .A1(n2756), .A2(n12882), .Y(n3189) );
  OR2X1_RVT U3135 ( .A1(n3191), .A2(n51), .Y(n3186) );
  AND2X1_RVT U3136 ( .A1(n2980), .A2(n2857), .Y(n3191) );
  OR2X1_RVT U3137 ( .A1(n2706), .A2(n3192), .Y(n2857) );
  OR2X1_RVT U3138 ( .A1(n12893), .A2(n12479), .Y(n3192) );
  AND4X1_RVT U3139 ( .A1(n2874), .A2(n3193), .A3(n3066), .A4(n3194), .Y(n3157)
         );
  AND4X1_RVT U3140 ( .A1(n3195), .A2(n3196), .A3(n3197), .A4(n3198), .Y(n3194)
         );
  OR2X1_RVT U3141 ( .A1(n2837), .A2(n2758), .Y(n3198) );
  OR2X1_RVT U3142 ( .A1(n2775), .A2(n2804), .Y(n3197) );
  OR2X1_RVT U3143 ( .A1(n12881), .A2(n3029), .Y(n3196) );
  OR2X1_RVT U3144 ( .A1(n2753), .A2(n2735), .Y(n3029) );
  OR2X1_RVT U3145 ( .A1(n12889), .A2(n2817), .Y(n2735) );
  OR2X1_RVT U3146 ( .A1(n12493), .A2(n2858), .Y(n3195) );
  OR2X1_RVT U3147 ( .A1(n2739), .A2(n2967), .Y(n2858) );
  OR2X1_RVT U3148 ( .A1(n12477), .A2(n2943), .Y(n2967) );
  AND2X1_RVT U3149 ( .A1(n3199), .A2(n3200), .Y(n3066) );
  OR2X1_RVT U3150 ( .A1(n3201), .A2(n2806), .Y(n3200) );
  OR2X1_RVT U3151 ( .A1(n12503), .A2(n51), .Y(n3201) );
  OR2X1_RVT U3152 ( .A1(n3202), .A2(n2689), .Y(n3199) );
  OR2X1_RVT U3153 ( .A1(n12880), .A2(n2806), .Y(n2689) );
  OR2X1_RVT U3154 ( .A1(n2703), .A2(n2753), .Y(n3202) );
  OR2X1_RVT U3155 ( .A1(n12485), .A2(n3072), .Y(n3193) );
  AND2X1_RVT U3156 ( .A1(n3203), .A2(n3204), .Y(n2874) );
  OR2X1_RVT U3157 ( .A1(n2757), .A2(n2795), .Y(n3204) );
  OR2X1_RVT U3158 ( .A1(n3205), .A2(n3206), .Y(n3203) );
  AND4X1_RVT U3159 ( .A1(n3207), .A2(n3208), .A3(n3209), .A4(n3210), .Y(n3156)
         );
  OR2X1_RVT U3160 ( .A1(n3211), .A2(n2943), .Y(n3210) );
  AND2X1_RVT U3161 ( .A1(n3212), .A2(n2952), .Y(n3211) );
  OR2X1_RVT U3162 ( .A1(n12491), .A2(n3168), .Y(n2952) );
  OR2X1_RVT U3163 ( .A1(n3213), .A2(n12886), .Y(n3209) );
  AND2X1_RVT U3164 ( .A1(n2880), .A2(n2845), .Y(n3213) );
  OR2X1_RVT U3165 ( .A1(n12880), .A2(n2821), .Y(n2845) );
  OR2X1_RVT U3166 ( .A1(n3214), .A2(n2900), .Y(n3208) );
  AND2X1_RVT U3167 ( .A1(n3215), .A2(n3216), .Y(n3214) );
  OR2X1_RVT U3168 ( .A1(n12480), .A2(n2759), .Y(n3216) );
  AND2X1_RVT U3169 ( .A1(n3217), .A2(n2797), .Y(n3215) );
  OR2X1_RVT U3170 ( .A1(n49), .A2(n2756), .Y(n3217) );
  OR2X1_RVT U3171 ( .A1(n3218), .A2(n2697), .Y(n3207) );
  AND2X1_RVT U3172 ( .A1(n3219), .A2(n3220), .Y(n3218) );
  NAND2X1_RVT U3173 ( .A1(n2682), .A2(n3060), .Y(n3220) );
  AND2X1_RVT U3174 ( .A1(n3221), .A2(n2910), .Y(n3219) );
  OR2X1_RVT U3175 ( .A1(n2843), .A2(n3168), .Y(n2910) );
  OR2X1_RVT U3176 ( .A1(n12500), .A2(n3222), .Y(n3221) );
  AND4X1_RVT U3177 ( .A1(n3223), .A2(n3224), .A3(n3225), .A4(n3226), .Y(n3155)
         );
  OR2X1_RVT U3178 ( .A1(n3227), .A2(n2720), .Y(n3226) );
  AND2X1_RVT U3179 ( .A1(n3228), .A2(n2861), .Y(n3227) );
  AND2X1_RVT U3180 ( .A1(n3229), .A2(n2883), .Y(n3228) );
  OR2X1_RVT U3181 ( .A1(n51), .A2(n3206), .Y(n2883) );
  OR2X1_RVT U3182 ( .A1(n12479), .A2(n2817), .Y(n3206) );
  OR2X1_RVT U3183 ( .A1(n3230), .A2(n12496), .Y(n3225) );
  AND2X1_RVT U3184 ( .A1(n3231), .A2(n3232), .Y(n3230) );
  OR2X1_RVT U3185 ( .A1(n3233), .A2(n12878), .Y(n3232) );
  AND2X1_RVT U3186 ( .A1(n3234), .A2(n3235), .Y(n3233) );
  OR2X1_RVT U3187 ( .A1(n12478), .A2(n3094), .Y(n3235) );
  OR2X1_RVT U3188 ( .A1(n12885), .A2(n2740), .Y(n3234) );
  AND2X1_RVT U3189 ( .A1(n3236), .A2(n3237), .Y(n3231) );
  OR2X1_RVT U3190 ( .A1(n2706), .A2(n3238), .Y(n3236) );
  OR2X1_RVT U3191 ( .A1(n3239), .A2(n2740), .Y(n3224) );
  AND4X1_RVT U3192 ( .A1(n3240), .A2(n3241), .A3(n3242), .A4(n2706), .Y(n3239)
         );
  OR2X1_RVT U3193 ( .A1(n12886), .A2(n2756), .Y(n3242) );
  OR2X1_RVT U3194 ( .A1(n12490), .A2(n2775), .Y(n3241) );
  OR2X1_RVT U3195 ( .A1(n2828), .A2(n2806), .Y(n3240) );
  OR2X1_RVT U3196 ( .A1(n3243), .A2(n2682), .Y(n3223) );
  AND4X1_RVT U3197 ( .A1(n3107), .A2(n3244), .A3(n2905), .A4(n2821), .Y(n3243)
         );
  OR2X1_RVT U3198 ( .A1(n2775), .A2(n3238), .Y(n2905) );
  OR2X1_RVT U3199 ( .A1(n2943), .A2(n3150), .Y(n3244) );
  OR2X1_RVT U3200 ( .A1(n12484), .A2(n2908), .Y(n3107) );
  AND4X1_RVT U3201 ( .A1(n3246), .A2(n3247), .A3(n3248), .A4(n3249), .Y(n3245)
         );
  AND4X1_RVT U3202 ( .A1(n3250), .A2(n3251), .A3(n3252), .A4(n3253), .Y(n3249)
         );
  AND4X1_RVT U3203 ( .A1(n3254), .A2(n3255), .A3(n3256), .A4(n3257), .Y(n3253)
         );
  OR2X1_RVT U3204 ( .A1(n12570), .A2(n3259), .Y(n3252) );
  OR2X1_RVT U3205 ( .A1(n3260), .A2(n3261), .Y(n3250) );
  OR2X1_RVT U3206 ( .A1(n12736), .A2(n3262), .Y(n3261) );
  AND4X1_RVT U3207 ( .A1(n3263), .A2(n3264), .A3(n3265), .A4(n3266), .Y(n3248)
         );
  OR2X1_RVT U3208 ( .A1(n3267), .A2(n12734), .Y(n3266) );
  AND2X1_RVT U3209 ( .A1(n3268), .A2(n3269), .Y(n3267) );
  AND2X1_RVT U3210 ( .A1(n3270), .A2(n3271), .Y(n3265) );
  OR2X1_RVT U3211 ( .A1(n3272), .A2(n256), .Y(n3271) );
  AND2X1_RVT U3212 ( .A1(n3273), .A2(n3274), .Y(n3272) );
  OR2X1_RVT U3213 ( .A1(n12561), .A2(n3276), .Y(n3274) );
  OR2X1_RVT U3214 ( .A1(n3262), .A2(n3277), .Y(n3273) );
  OR2X1_RVT U3215 ( .A1(n3278), .A2(n12567), .Y(n3270) );
  AND2X1_RVT U3216 ( .A1(n3280), .A2(n3281), .Y(n3278) );
  OR2X1_RVT U3217 ( .A1(n3282), .A2(n3283), .Y(n3264) );
  AND2X1_RVT U3218 ( .A1(n3284), .A2(n3285), .Y(n3282) );
  OR2X1_RVT U3219 ( .A1(n12562), .A2(n3286), .Y(n3285) );
  AND2X1_RVT U3220 ( .A1(n3287), .A2(n3288), .Y(n3284) );
  AND2X1_RVT U3221 ( .A1(n3289), .A2(n3290), .Y(n3263) );
  OR2X1_RVT U3222 ( .A1(n3291), .A2(n12544), .Y(n3290) );
  AND2X1_RVT U3223 ( .A1(n3293), .A2(n3294), .Y(n3291) );
  OR2X1_RVT U3224 ( .A1(n3295), .A2(n3296), .Y(n3294) );
  OR2X1_RVT U3225 ( .A1(n12553), .A2(n12548), .Y(n3296) );
  OR2X1_RVT U3226 ( .A1(n3299), .A2(n3300), .Y(n3289) );
  AND2X1_RVT U3227 ( .A1(n3301), .A2(n3302), .Y(n3299) );
  AND2X1_RVT U3228 ( .A1(n3303), .A2(n3304), .Y(n3301) );
  AND4X1_RVT U3229 ( .A1(n3305), .A2(n3306), .A3(n3307), .A4(n3308), .Y(n3247)
         );
  AND4X1_RVT U3230 ( .A1(n3309), .A2(n3310), .A3(n3311), .A4(n3312), .Y(n3308)
         );
  OR2X1_RVT U3231 ( .A1(n3313), .A2(n12573), .Y(n3312) );
  AND4X1_RVT U3232 ( .A1(n3315), .A2(n3316), .A3(n3317), .A4(n3318), .Y(n3313)
         );
  OR2X1_RVT U3233 ( .A1(n3319), .A2(n3286), .Y(n3318) );
  OR2X1_RVT U3234 ( .A1(n3320), .A2(n12559), .Y(n3317) );
  OR2X1_RVT U3235 ( .A1(n3322), .A2(n12550), .Y(n3311) );
  AND4X1_RVT U3236 ( .A1(n3323), .A2(n3324), .A3(n3325), .A4(n3326), .Y(n3322)
         );
  OR2X1_RVT U3237 ( .A1(n3327), .A2(n3328), .Y(n3326) );
  OR2X1_RVT U3238 ( .A1(n12567), .A2(n12562), .Y(n3328) );
  AND2X1_RVT U3239 ( .A1(n3329), .A2(n3330), .Y(n3325) );
  OR2X1_RVT U3240 ( .A1(n12738), .A2(n3331), .Y(n3324) );
  OR2X1_RVT U3241 ( .A1(n3332), .A2(n3333), .Y(n3323) );
  AND2X1_RVT U3242 ( .A1(n3334), .A2(n3335), .Y(n3332) );
  OR2X1_RVT U3243 ( .A1(n12567), .A2(n3336), .Y(n3335) );
  OR2X1_RVT U3244 ( .A1(n3269), .A2(n3337), .Y(n3310) );
  OR2X1_RVT U3245 ( .A1(n3336), .A2(n3338), .Y(n3309) );
  OR2X1_RVT U3246 ( .A1(n3339), .A2(n3340), .Y(n3307) );
  OR2X1_RVT U3247 ( .A1(n3341), .A2(n3334), .Y(n3306) );
  OR2X1_RVT U3248 ( .A1(n3342), .A2(n3343), .Y(n3305) );
  AND4X1_RVT U3249 ( .A1(n3344), .A2(n3345), .A3(n3346), .A4(n3347), .Y(n3246)
         );
  AND2X1_RVT U3250 ( .A1(n3348), .A2(n3349), .Y(n3347) );
  OR2X1_RVT U3251 ( .A1(n3333), .A2(n3350), .Y(n3349) );
  AND2X1_RVT U3252 ( .A1(n3351), .A2(n3352), .Y(n3348) );
  OR2X1_RVT U3253 ( .A1(n3353), .A2(n3276), .Y(n3352) );
  OR2X1_RVT U3254 ( .A1(n3277), .A2(n3354), .Y(n3351) );
  OR2X1_RVT U3255 ( .A1(n254), .A2(n3355), .Y(n3346) );
  OR2X1_RVT U3256 ( .A1(n3356), .A2(n12557), .Y(n3345) );
  OR2X1_RVT U3257 ( .A1(n12560), .A2(n3358), .Y(n3344) );
  AND4X1_RVT U3258 ( .A1(n3360), .A2(n3361), .A3(n3362), .A4(n3363), .Y(n3359)
         );
  AND4X1_RVT U3259 ( .A1(n3364), .A2(n3255), .A3(n3365), .A4(n3366), .Y(n3363)
         );
  AND4X1_RVT U3260 ( .A1(n3367), .A2(n3368), .A3(n3369), .A4(n3370), .Y(n3366)
         );
  OR2X1_RVT U3261 ( .A1(n3276), .A2(n3371), .Y(n3370) );
  OR2X1_RVT U3262 ( .A1(n3372), .A2(n12572), .Y(n3371) );
  OR2X1_RVT U3263 ( .A1(n3277), .A2(n3373), .Y(n3369) );
  OR2X1_RVT U3264 ( .A1(n254), .A2(n12556), .Y(n3373) );
  OR2X1_RVT U3265 ( .A1(n3374), .A2(n3320), .Y(n3368) );
  AND2X1_RVT U3266 ( .A1(n3331), .A2(n3375), .Y(n3374) );
  OR2X1_RVT U3267 ( .A1(n3376), .A2(n3377), .Y(n3367) );
  AND2X1_RVT U3268 ( .A1(n3378), .A2(n3379), .Y(n3376) );
  AND2X1_RVT U3269 ( .A1(n3380), .A2(n3381), .Y(n3365) );
  OR2X1_RVT U3270 ( .A1(n3327), .A2(n3382), .Y(n3381) );
  OR2X1_RVT U3271 ( .A1(n3383), .A2(n12736), .Y(n3382) );
  OR2X1_RVT U3272 ( .A1(n3384), .A2(n3385), .Y(n3380) );
  OR2X1_RVT U3273 ( .A1(n3386), .A2(n12561), .Y(n3385) );
  OR2X1_RVT U3274 ( .A1(n3262), .A2(n3387), .Y(n3255) );
  AND4X1_RVT U3275 ( .A1(n3388), .A2(n3389), .A3(n3390), .A4(n3391), .Y(n3362)
         );
  AND4X1_RVT U3276 ( .A1(n3392), .A2(n3393), .A3(n3394), .A4(n3395), .Y(n3391)
         );
  OR2X1_RVT U3277 ( .A1(n3396), .A2(n12575), .Y(n3395) );
  AND2X1_RVT U3278 ( .A1(n3398), .A2(n3399), .Y(n3396) );
  OR2X1_RVT U3279 ( .A1(n12544), .A2(n3277), .Y(n3399) );
  OR2X1_RVT U3280 ( .A1(n3400), .A2(n3279), .Y(n3394) );
  AND2X1_RVT U3281 ( .A1(n3401), .A2(n3402), .Y(n3400) );
  OR2X1_RVT U3282 ( .A1(n3403), .A2(n12735), .Y(n3393) );
  AND2X1_RVT U3283 ( .A1(n3404), .A2(n3405), .Y(n3403) );
  OR2X1_RVT U3284 ( .A1(n3406), .A2(n3355), .Y(n3405) );
  AND2X1_RVT U3285 ( .A1(n12575), .A2(n12559), .Y(n3406) );
  OR2X1_RVT U3286 ( .A1(n3407), .A2(n12545), .Y(n3392) );
  AND2X1_RVT U3287 ( .A1(n3409), .A2(n3410), .Y(n3407) );
  OR2X1_RVT U3288 ( .A1(n3411), .A2(n12551), .Y(n3390) );
  AND2X1_RVT U3289 ( .A1(n3412), .A2(n3413), .Y(n3411) );
  OR2X1_RVT U3290 ( .A1(n12559), .A2(n3414), .Y(n3413) );
  AND2X1_RVT U3291 ( .A1(n3415), .A2(n3416), .Y(n3412) );
  OR2X1_RVT U3292 ( .A1(n3417), .A2(n3418), .Y(n3415) );
  OR2X1_RVT U3293 ( .A1(n3262), .A2(n3333), .Y(n3418) );
  OR2X1_RVT U3294 ( .A1(n3419), .A2(n12732), .Y(n3389) );
  AND2X1_RVT U3295 ( .A1(n3420), .A2(n3421), .Y(n3419) );
  OR2X1_RVT U3296 ( .A1(n3422), .A2(n3423), .Y(n3388) );
  AND2X1_RVT U3297 ( .A1(n3424), .A2(n3425), .Y(n3422) );
  AND2X1_RVT U3298 ( .A1(n3426), .A2(n3427), .Y(n3424) );
  OR2X1_RVT U3299 ( .A1(n256), .A2(n3355), .Y(n3427) );
  OR2X1_RVT U3300 ( .A1(n12569), .A2(n3320), .Y(n3426) );
  AND4X1_RVT U3301 ( .A1(n3428), .A2(n3429), .A3(n3430), .A4(n3431), .Y(n3361)
         );
  AND4X1_RVT U3302 ( .A1(n3432), .A2(n3433), .A3(n3434), .A4(n3435), .Y(n3431)
         );
  OR2X1_RVT U3303 ( .A1(n3355), .A2(n3354), .Y(n3435) );
  OR2X1_RVT U3304 ( .A1(n3286), .A2(n3436), .Y(n3434) );
  OR2X1_RVT U3305 ( .A1(n3319), .A2(n3437), .Y(n3433) );
  OR2X1_RVT U3306 ( .A1(n3262), .A2(n3438), .Y(n3432) );
  AND2X1_RVT U3307 ( .A1(n3439), .A2(n3440), .Y(n3430) );
  OR2X1_RVT U3308 ( .A1(n12570), .A2(n3441), .Y(n3440) );
  OR2X1_RVT U3309 ( .A1(n12549), .A2(n3338), .Y(n3439) );
  OR2X1_RVT U3310 ( .A1(n3442), .A2(n3297), .Y(n3429) );
  AND4X1_RVT U3311 ( .A1(n3443), .A2(n3444), .A3(n3445), .A4(n3446), .Y(n3442)
         );
  OR2X1_RVT U3312 ( .A1(n3447), .A2(n3262), .Y(n3445) );
  OR2X1_RVT U3313 ( .A1(n12724), .A2(n3448), .Y(n3444) );
  OR2X1_RVT U3314 ( .A1(n3449), .A2(n12732), .Y(n3443) );
  AND2X1_RVT U3315 ( .A1(n3340), .A2(n3450), .Y(n3449) );
  OR2X1_RVT U3316 ( .A1(n3342), .A2(n3451), .Y(n3428) );
  AND4X1_RVT U3317 ( .A1(n3452), .A2(n3453), .A3(n3454), .A4(n3455), .Y(n3360)
         );
  AND4X1_RVT U3318 ( .A1(n3456), .A2(n3457), .A3(n3458), .A4(n3459), .Y(n3455)
         );
  OR2X1_RVT U3319 ( .A1(n12728), .A2(n3460), .Y(n3459) );
  OR2X1_RVT U3320 ( .A1(n12729), .A2(n3461), .Y(n3458) );
  OR2X1_RVT U3321 ( .A1(n12726), .A2(n3462), .Y(n3457) );
  OR2X1_RVT U3322 ( .A1(n12543), .A2(n3463), .Y(n3456) );
  OR2X1_RVT U3323 ( .A1(n3464), .A2(n12550), .Y(n3453) );
  AND4X1_RVT U3324 ( .A1(n3466), .A2(n3467), .A3(n3468), .A4(n3469), .Y(n3465)
         );
  AND4X1_RVT U3325 ( .A1(n3470), .A2(n3471), .A3(n3472), .A4(n3473), .Y(n3469)
         );
  AND4X1_RVT U3326 ( .A1(n3474), .A2(n3251), .A3(n3421), .A4(n3475), .Y(n3473)
         );
  OR2X1_RVT U3327 ( .A1(n3476), .A2(n12723), .Y(n3251) );
  AND2X1_RVT U3328 ( .A1(n3477), .A2(n3478), .Y(n3476) );
  OR2X1_RVT U3329 ( .A1(n3295), .A2(n3479), .Y(n3478) );
  OR2X1_RVT U3330 ( .A1(n3480), .A2(n3377), .Y(n3477) );
  OR2X1_RVT U3331 ( .A1(n3481), .A2(n3336), .Y(n3474) );
  AND2X1_RVT U3332 ( .A1(n3482), .A2(n3483), .Y(n3481) );
  OR2X1_RVT U3333 ( .A1(n12728), .A2(n3320), .Y(n3483) );
  OR2X1_RVT U3334 ( .A1(n3484), .A2(n3279), .Y(n3472) );
  AND2X1_RVT U3335 ( .A1(n3485), .A2(n3486), .Y(n3484) );
  OR2X1_RVT U3336 ( .A1(n3487), .A2(n12734), .Y(n3486) );
  AND2X1_RVT U3337 ( .A1(n3327), .A2(n3488), .Y(n3487) );
  OR2X1_RVT U3338 ( .A1(n3489), .A2(n12570), .Y(n3471) );
  AND2X1_RVT U3339 ( .A1(n3490), .A2(n3491), .Y(n3489) );
  OR2X1_RVT U3340 ( .A1(n3320), .A2(n3286), .Y(n3491) );
  OR2X1_RVT U3341 ( .A1(n3492), .A2(n12553), .Y(n3470) );
  AND2X1_RVT U3342 ( .A1(n3404), .A2(n3493), .Y(n3492) );
  OR2X1_RVT U3343 ( .A1(n3333), .A2(n3494), .Y(n3404) );
  AND4X1_RVT U3344 ( .A1(n3495), .A2(n3496), .A3(n3497), .A4(n3498), .Y(n3468)
         );
  OR2X1_RVT U3345 ( .A1(n3499), .A2(n12560), .Y(n3498) );
  AND2X1_RVT U3346 ( .A1(n3500), .A2(n3501), .Y(n3499) );
  OR2X1_RVT U3347 ( .A1(n3377), .A2(n3277), .Y(n3501) );
  AND2X1_RVT U3348 ( .A1(n3502), .A2(n3503), .Y(n3500) );
  OR2X1_RVT U3349 ( .A1(n3417), .A2(n3479), .Y(n3502) );
  AND2X1_RVT U3350 ( .A1(n3504), .A2(n3505), .Y(n3497) );
  OR2X1_RVT U3351 ( .A1(n3506), .A2(n3408), .Y(n3505) );
  AND2X1_RVT U3352 ( .A1(n3507), .A2(n3316), .Y(n3506) );
  OR2X1_RVT U3353 ( .A1(n3262), .A2(n3377), .Y(n3316) );
  OR2X1_RVT U3354 ( .A1(n3508), .A2(n256), .Y(n3504) );
  AND2X1_RVT U3355 ( .A1(n3509), .A2(n3510), .Y(n3508) );
  OR2X1_RVT U3356 ( .A1(n3511), .A2(n12562), .Y(n3510) );
  AND2X1_RVT U3357 ( .A1(n3512), .A2(n3513), .Y(n3511) );
  OR2X1_RVT U3358 ( .A1(n12557), .A2(n3327), .Y(n3513) );
  OR2X1_RVT U3359 ( .A1(n12738), .A2(n12559), .Y(n3512) );
  AND2X1_RVT U3360 ( .A1(n3378), .A2(n3488), .Y(n3509) );
  OR2X1_RVT U3361 ( .A1(n3408), .A2(n3514), .Y(n3378) );
  OR2X1_RVT U3362 ( .A1(n12733), .A2(n12729), .Y(n3514) );
  OR2X1_RVT U3363 ( .A1(n3515), .A2(n3397), .Y(n3496) );
  AND4X1_RVT U3364 ( .A1(n3356), .A2(n3516), .A3(n3517), .A4(n3518), .Y(n3515)
         );
  OR2X1_RVT U3365 ( .A1(n12561), .A2(n3377), .Y(n3518) );
  AND2X1_RVT U3366 ( .A1(n3519), .A2(n3520), .Y(n3517) );
  OR2X1_RVT U3367 ( .A1(n12738), .A2(n12570), .Y(n3516) );
  AND2X1_RVT U3368 ( .A1(n3521), .A2(n3522), .Y(n3356) );
  OR2X1_RVT U3369 ( .A1(n3523), .A2(n254), .Y(n3522) );
  OR2X1_RVT U3370 ( .A1(n3320), .A2(n12723), .Y(n3521) );
  AND2X1_RVT U3371 ( .A1(n3524), .A2(n3525), .Y(n3495) );
  OR2X1_RVT U3372 ( .A1(n3526), .A2(n12725), .Y(n3525) );
  AND2X1_RVT U3373 ( .A1(n3527), .A2(n3528), .Y(n3526) );
  OR2X1_RVT U3374 ( .A1(n3529), .A2(n12564), .Y(n3528) );
  AND2X1_RVT U3375 ( .A1(n3530), .A2(n3531), .Y(n3529) );
  AND2X1_RVT U3376 ( .A1(n3532), .A2(n3533), .Y(n3527) );
  OR2X1_RVT U3377 ( .A1(n3534), .A2(n12573), .Y(n3524) );
  AND4X1_RVT U3378 ( .A1(n3535), .A2(n3536), .A3(n3537), .A4(n3538), .Y(n3534)
         );
  OR2X1_RVT U3379 ( .A1(n12737), .A2(n3539), .Y(n3537) );
  OR2X1_RVT U3380 ( .A1(n254), .A2(n3334), .Y(n3536) );
  OR2X1_RVT U3381 ( .A1(n3423), .A2(n3377), .Y(n3535) );
  AND4X1_RVT U3382 ( .A1(n3540), .A2(n3541), .A3(n3542), .A4(n3543), .Y(n3467)
         );
  AND2X1_RVT U3383 ( .A1(n3544), .A2(n3387), .Y(n3543) );
  OR2X1_RVT U3384 ( .A1(n12548), .A2(n3353), .Y(n3387) );
  AND2X1_RVT U3385 ( .A1(n3545), .A2(n3546), .Y(n3544) );
  OR2X1_RVT U3386 ( .A1(n3547), .A2(n3302), .Y(n3546) );
  OR2X1_RVT U3387 ( .A1(n3354), .A2(n3414), .Y(n3545) );
  OR2X1_RVT U3388 ( .A1(n254), .A2(n3548), .Y(n3542) );
  OR2X1_RVT U3389 ( .A1(n12736), .A2(n3549), .Y(n3541) );
  OR2X1_RVT U3390 ( .A1(n3423), .A2(n3550), .Y(n3540) );
  AND4X1_RVT U3391 ( .A1(n3551), .A2(n3552), .A3(n3553), .A4(n3554), .Y(n3466)
         );
  AND2X1_RVT U3392 ( .A1(n3555), .A2(n3556), .Y(n3554) );
  OR2X1_RVT U3393 ( .A1(n12543), .A2(n3557), .Y(n3556) );
  AND2X1_RVT U3394 ( .A1(n3558), .A2(n3559), .Y(n3555) );
  OR2X1_RVT U3395 ( .A1(n3319), .A2(n3329), .Y(n3559) );
  OR2X1_RVT U3396 ( .A1(n12564), .A2(n3379), .Y(n3329) );
  OR2X1_RVT U3397 ( .A1(n12550), .A2(n3560), .Y(n3558) );
  OR2X1_RVT U3398 ( .A1(n3300), .A2(n3293), .Y(n3553) );
  OR2X1_RVT U3399 ( .A1(n3386), .A2(n3561), .Y(n3293) );
  OR2X1_RVT U3400 ( .A1(n12732), .A2(n3562), .Y(n3552) );
  OR2X1_RVT U3401 ( .A1(n12562), .A2(n3420), .Y(n3551) );
  OR2X1_RVT U3402 ( .A1(n12723), .A2(n3482), .Y(n3420) );
  AND4X1_RVT U3403 ( .A1(n3564), .A2(n3565), .A3(n3566), .A4(n3567), .Y(n3563)
         );
  AND4X1_RVT U3404 ( .A1(n3568), .A2(n3569), .A3(n3570), .A4(n3571), .Y(n3567)
         );
  OR2X1_RVT U3405 ( .A1(n264), .A2(n3572), .Y(n3571) );
  OR2X1_RVT U3406 ( .A1(n3573), .A2(n12575), .Y(n3572) );
  AND2X1_RVT U3407 ( .A1(n12564), .A2(n3339), .Y(n3573) );
  AND2X1_RVT U3408 ( .A1(n3254), .A2(n3574), .Y(n3570) );
  OR2X1_RVT U3409 ( .A1(n12553), .A2(n3575), .Y(n3254) );
  OR2X1_RVT U3410 ( .A1(n264), .A2(n3333), .Y(n3575) );
  OR2X1_RVT U3411 ( .A1(n3576), .A2(n3262), .Y(n3569) );
  AND2X1_RVT U3412 ( .A1(n3577), .A2(n3578), .Y(n3576) );
  AND2X1_RVT U3413 ( .A1(n3579), .A2(n3580), .Y(n3568) );
  OR2X1_RVT U3414 ( .A1(n3581), .A2(n3582), .Y(n3580) );
  AND2X1_RVT U3415 ( .A1(n3583), .A2(n3343), .Y(n3581) );
  OR2X1_RVT U3416 ( .A1(n3584), .A2(n3334), .Y(n3579) );
  AND2X1_RVT U3417 ( .A1(n3519), .A2(n3353), .Y(n3584) );
  OR2X1_RVT U3418 ( .A1(n12551), .A2(n3585), .Y(n3519) );
  OR2X1_RVT U3419 ( .A1(n12738), .A2(n12561), .Y(n3585) );
  AND4X1_RVT U3420 ( .A1(n3586), .A2(n3587), .A3(n3588), .A4(n3589), .Y(n3566)
         );
  OR2X1_RVT U3421 ( .A1(n3590), .A2(n12728), .Y(n3589) );
  AND2X1_RVT U3422 ( .A1(n3402), .A2(n3591), .Y(n3590) );
  OR2X1_RVT U3423 ( .A1(n12736), .A2(n3447), .Y(n3402) );
  AND2X1_RVT U3424 ( .A1(n3592), .A2(n3593), .Y(n3588) );
  OR2X1_RVT U3425 ( .A1(n3594), .A2(n12726), .Y(n3593) );
  AND2X1_RVT U3426 ( .A1(n3595), .A2(n3596), .Y(n3594) );
  OR2X1_RVT U3427 ( .A1(n3297), .A2(n3539), .Y(n3596) );
  OR2X1_RVT U3428 ( .A1(n3597), .A2(n12724), .Y(n3592) );
  AND2X1_RVT U3429 ( .A1(n3598), .A2(n3599), .Y(n3597) );
  OR2X1_RVT U3430 ( .A1(n3600), .A2(n12564), .Y(n3587) );
  AND2X1_RVT U3431 ( .A1(n3601), .A2(n3602), .Y(n3600) );
  AND2X1_RVT U3432 ( .A1(n3603), .A2(n3604), .Y(n3601) );
  AND2X1_RVT U3433 ( .A1(n3605), .A2(n3606), .Y(n3586) );
  OR2X1_RVT U3434 ( .A1(n3607), .A2(n3523), .Y(n3606) );
  AND2X1_RVT U3435 ( .A1(n3608), .A2(n3354), .Y(n3607) );
  AND2X1_RVT U3436 ( .A1(n3609), .A2(n3610), .Y(n3608) );
  OR2X1_RVT U3437 ( .A1(n3611), .A2(n12567), .Y(n3605) );
  AND2X1_RVT U3438 ( .A1(n3612), .A2(n3613), .Y(n3611) );
  OR2X1_RVT U3439 ( .A1(n12735), .A2(n12569), .Y(n3613) );
  AND2X1_RVT U3440 ( .A1(n3343), .A2(n3614), .Y(n3612) );
  AND4X1_RVT U3441 ( .A1(n3615), .A2(n3616), .A3(n3617), .A4(n3618), .Y(n3565)
         );
  AND2X1_RVT U3442 ( .A1(n3619), .A2(n3620), .Y(n3618) );
  OR2X1_RVT U3443 ( .A1(n3336), .A2(n3410), .Y(n3620) );
  OR2X1_RVT U3444 ( .A1(n12730), .A2(n3343), .Y(n3410) );
  AND2X1_RVT U3445 ( .A1(n3621), .A2(n3622), .Y(n3619) );
  OR2X1_RVT U3446 ( .A1(n3488), .A2(n3302), .Y(n3622) );
  OR2X1_RVT U3447 ( .A1(n12737), .A2(n12560), .Y(n3302) );
  OR2X1_RVT U3448 ( .A1(n3386), .A2(n3436), .Y(n3621) );
  OR2X1_RVT U3449 ( .A1(n12725), .A2(n3623), .Y(n3436) );
  OR2X1_RVT U3450 ( .A1(n3624), .A2(n12543), .Y(n3617) );
  AND4X1_RVT U3451 ( .A1(n3625), .A2(n3626), .A3(n3627), .A4(n3628), .Y(n3624)
         );
  OR2X1_RVT U3452 ( .A1(n3561), .A2(n3334), .Y(n3627) );
  OR2X1_RVT U3453 ( .A1(n3629), .A2(n3331), .Y(n3626) );
  OR2X1_RVT U3454 ( .A1(n12734), .A2(n3286), .Y(n3625) );
  OR2X1_RVT U3455 ( .A1(n3630), .A2(n12544), .Y(n3616) );
  AND2X1_RVT U3456 ( .A1(n3631), .A2(n3632), .Y(n3630) );
  OR2X1_RVT U3457 ( .A1(n3561), .A2(n3286), .Y(n3632) );
  AND2X1_RVT U3458 ( .A1(n3633), .A2(n3562), .Y(n3631) );
  OR2X1_RVT U3459 ( .A1(n3334), .A2(n3634), .Y(n3562) );
  OR2X1_RVT U3460 ( .A1(n12725), .A2(n12737), .Y(n3634) );
  OR2X1_RVT U3461 ( .A1(n3635), .A2(n12551), .Y(n3615) );
  AND4X1_RVT U3462 ( .A1(n3636), .A2(n3549), .A3(n3358), .A4(n3330), .Y(n3635)
         );
  OR2X1_RVT U3463 ( .A1(n3355), .A2(n3637), .Y(n3330) );
  OR2X1_RVT U3464 ( .A1(n12727), .A2(n3292), .Y(n3637) );
  OR2X1_RVT U3465 ( .A1(n3417), .A2(n3451), .Y(n3358) );
  OR2X1_RVT U3466 ( .A1(n3336), .A2(n3638), .Y(n3549) );
  OR2X1_RVT U3467 ( .A1(n12575), .A2(n12544), .Y(n3638) );
  OR2X1_RVT U3468 ( .A1(n3295), .A2(n3639), .Y(n3636) );
  OR2X1_RVT U3469 ( .A1(n3640), .A2(n12549), .Y(n3639) );
  AND4X1_RVT U3470 ( .A1(n3641), .A2(n3642), .A3(n3643), .A4(n3644), .Y(n3564)
         );
  AND2X1_RVT U3471 ( .A1(n3645), .A2(n3646), .Y(n3644) );
  AND2X1_RVT U3472 ( .A1(n3647), .A2(n3648), .Y(n3645) );
  OR2X1_RVT U3473 ( .A1(n3327), .A2(n3602), .Y(n3648) );
  OR2X1_RVT U3474 ( .A1(n3339), .A2(n3649), .Y(n3602) );
  OR2X1_RVT U3475 ( .A1(n12726), .A2(n12728), .Y(n3649) );
  OR2X1_RVT U3476 ( .A1(n12733), .A2(n3650), .Y(n3647) );
  OR2X1_RVT U3477 ( .A1(n12560), .A2(n3651), .Y(n3643) );
  OR2X1_RVT U3478 ( .A1(n12736), .A2(n3652), .Y(n3642) );
  OR2X1_RVT U3479 ( .A1(n3339), .A2(n3653), .Y(n3641) );
  AND4X1_RVT U3480 ( .A1(n3655), .A2(n3656), .A3(n3657), .A4(n3658), .Y(n3654)
         );
  AND4X1_RVT U3481 ( .A1(n3659), .A2(n3660), .A3(n3661), .A4(n3662), .Y(n3658)
         );
  AND4X1_RVT U3482 ( .A1(n3663), .A2(n3664), .A3(n3256), .A4(n3665), .Y(n3662)
         );
  OR2X1_RVT U3483 ( .A1(n3397), .A2(n3666), .Y(n3256) );
  OR2X1_RVT U3484 ( .A1(n3488), .A2(n256), .Y(n3666) );
  OR2X1_RVT U3485 ( .A1(n3260), .A2(n3667), .Y(n3664) );
  OR2X1_RVT U3486 ( .A1(n12731), .A2(n12734), .Y(n3667) );
  OR2X1_RVT U3487 ( .A1(n3523), .A2(n3668), .Y(n3663) );
  OR2X1_RVT U3488 ( .A1(n3669), .A2(n3297), .Y(n3668) );
  AND2X1_RVT U3489 ( .A1(n12564), .A2(n3397), .Y(n3669) );
  OR2X1_RVT U3490 ( .A1(n3670), .A2(n12570), .Y(n3661) );
  AND2X1_RVT U3491 ( .A1(n3538), .A2(n3610), .Y(n3670) );
  OR2X1_RVT U3492 ( .A1(n256), .A2(n3671), .Y(n3610) );
  OR2X1_RVT U3493 ( .A1(n12543), .A2(n12730), .Y(n3671) );
  OR2X1_RVT U3494 ( .A1(n3327), .A2(n3672), .Y(n3538) );
  OR2X1_RVT U3495 ( .A1(n12728), .A2(n3319), .Y(n3672) );
  OR2X1_RVT U3496 ( .A1(n3673), .A2(n3277), .Y(n3660) );
  AND2X1_RVT U3497 ( .A1(n3674), .A2(n3482), .Y(n3673) );
  OR2X1_RVT U3498 ( .A1(n3383), .A2(n3377), .Y(n3659) );
  AND4X1_RVT U3499 ( .A1(n3675), .A2(n3676), .A3(n3677), .A4(n3678), .Y(n3657)
         );
  AND2X1_RVT U3500 ( .A1(n3679), .A2(n3680), .Y(n3678) );
  OR2X1_RVT U3501 ( .A1(n3681), .A2(n12564), .Y(n3680) );
  AND2X1_RVT U3502 ( .A1(n3682), .A2(n3350), .Y(n3681) );
  AND2X1_RVT U3503 ( .A1(n3683), .A2(n3684), .Y(n3679) );
  OR2X1_RVT U3504 ( .A1(n3685), .A2(n3333), .Y(n3684) );
  AND2X1_RVT U3505 ( .A1(n3304), .A2(n3276), .Y(n3685) );
  OR2X1_RVT U3506 ( .A1(n12736), .A2(n3375), .Y(n3304) );
  OR2X1_RVT U3507 ( .A1(n3686), .A2(n3386), .Y(n3683) );
  AND2X1_RVT U3508 ( .A1(n3578), .A2(n3687), .Y(n3686) );
  OR2X1_RVT U3509 ( .A1(n12737), .A2(n3414), .Y(n3578) );
  OR2X1_RVT U3510 ( .A1(n3688), .A2(n12728), .Y(n3677) );
  AND2X1_RVT U3511 ( .A1(n3281), .A2(n3689), .Y(n3688) );
  OR2X1_RVT U3512 ( .A1(n3417), .A2(n3341), .Y(n3689) );
  OR2X1_RVT U3513 ( .A1(n3320), .A2(n3523), .Y(n3281) );
  OR2X1_RVT U3514 ( .A1(n3690), .A2(n254), .Y(n3676) );
  AND2X1_RVT U3515 ( .A1(n3331), .A2(n3691), .Y(n3690) );
  OR2X1_RVT U3516 ( .A1(n3692), .A2(n12548), .Y(n3691) );
  AND2X1_RVT U3517 ( .A1(n3693), .A2(n3694), .Y(n3692) );
  OR2X1_RVT U3518 ( .A1(n12729), .A2(n3314), .Y(n3694) );
  OR2X1_RVT U3519 ( .A1(n12575), .A2(n3417), .Y(n3331) );
  OR2X1_RVT U3520 ( .A1(n3695), .A2(n3401), .Y(n3675) );
  AND2X1_RVT U3521 ( .A1(n3334), .A2(n3379), .Y(n3695) );
  OR2X1_RVT U3522 ( .A1(n12725), .A2(n3262), .Y(n3379) );
  AND4X1_RVT U3523 ( .A1(n3696), .A2(n3697), .A3(n3698), .A4(n3699), .Y(n3656)
         );
  AND4X1_RVT U3524 ( .A1(n3700), .A2(n3701), .A3(n3702), .A4(n3703), .Y(n3699)
         );
  OR2X1_RVT U3525 ( .A1(n3704), .A2(n12736), .Y(n3703) );
  AND2X1_RVT U3526 ( .A1(n3437), .A2(n3705), .Y(n3704) );
  OR2X1_RVT U3527 ( .A1(n12572), .A2(n3286), .Y(n3705) );
  OR2X1_RVT U3528 ( .A1(n3706), .A2(n3279), .Y(n3702) );
  AND2X1_RVT U3529 ( .A1(n3707), .A2(n3708), .Y(n3706) );
  OR2X1_RVT U3530 ( .A1(n3709), .A2(n3314), .Y(n3708) );
  AND2X1_RVT U3531 ( .A1(n3339), .A2(n3327), .Y(n3709) );
  AND2X1_RVT U3532 ( .A1(n3341), .A2(n3583), .Y(n3707) );
  OR2X1_RVT U3533 ( .A1(n12573), .A2(n3479), .Y(n3583) );
  OR2X1_RVT U3534 ( .A1(n3710), .A2(n12562), .Y(n3701) );
  AND2X1_RVT U3535 ( .A1(n3711), .A2(n3712), .Y(n3710) );
  OR2X1_RVT U3536 ( .A1(n3327), .A2(n3713), .Y(n3712) );
  AND2X1_RVT U3537 ( .A1(n3409), .A2(n3603), .Y(n3711) );
  OR2X1_RVT U3538 ( .A1(n3319), .A2(n3494), .Y(n3603) );
  OR2X1_RVT U3539 ( .A1(n3292), .A2(n3714), .Y(n3409) );
  OR2X1_RVT U3540 ( .A1(n3715), .A2(n3262), .Y(n3700) );
  AND4X1_RVT U3541 ( .A1(n3716), .A2(n3717), .A3(n3718), .A4(n3651), .Y(n3715)
         );
  OR2X1_RVT U3542 ( .A1(n3355), .A2(n3719), .Y(n3651) );
  OR2X1_RVT U3543 ( .A1(n12543), .A2(n3319), .Y(n3719) );
  OR2X1_RVT U3544 ( .A1(n12733), .A2(n3561), .Y(n3717) );
  OR2X1_RVT U3545 ( .A1(n3320), .A2(n3417), .Y(n3716) );
  OR2X1_RVT U3546 ( .A1(n3488), .A2(n3530), .Y(n3698) );
  OR2X1_RVT U3547 ( .A1(n3720), .A2(n12546), .Y(n3697) );
  AND4X1_RVT U3548 ( .A1(n3721), .A2(n3722), .A3(n3364), .A4(n3462), .Y(n3720)
         );
  OR2X1_RVT U3549 ( .A1(n3286), .A2(n3451), .Y(n3462) );
  OR2X1_RVT U3550 ( .A1(n12733), .A2(n254), .Y(n3451) );
  OR2X1_RVT U3551 ( .A1(n3279), .A2(n3343), .Y(n3364) );
  OR2X1_RVT U3552 ( .A1(n12725), .A2(n3714), .Y(n3696) );
  AND4X1_RVT U3553 ( .A1(n3723), .A2(n3724), .A3(n3725), .A4(n3726), .Y(n3655)
         );
  OR2X1_RVT U3554 ( .A1(n12551), .A2(n3727), .Y(n3726) );
  AND2X1_RVT U3555 ( .A1(n3728), .A2(n3729), .Y(n3725) );
  OR2X1_RVT U3556 ( .A1(n12572), .A2(n3482), .Y(n3729) );
  OR2X1_RVT U3557 ( .A1(n3269), .A2(n3343), .Y(n3728) );
  OR2X1_RVT U3558 ( .A1(n256), .A2(n3300), .Y(n3343) );
  OR2X1_RVT U3559 ( .A1(n12575), .A2(n3461), .Y(n3724) );
  OR2X1_RVT U3560 ( .A1(n3336), .A2(n3730), .Y(n3461) );
  AND2X1_RVT U3561 ( .A1(n3731), .A2(n3732), .Y(n3723) );
  OR2X1_RVT U3562 ( .A1(n12544), .A2(n3733), .Y(n3732) );
  OR2X1_RVT U3563 ( .A1(n3339), .A2(n3288), .Y(n3731) );
  OR2X1_RVT U3564 ( .A1(n3262), .A2(n3547), .Y(n3288) );
  AND4X1_RVT U3565 ( .A1(n3735), .A2(n3736), .A3(n3737), .A4(n3738), .Y(n3734)
         );
  AND4X1_RVT U3566 ( .A1(n3739), .A2(n3740), .A3(n3741), .A4(n3742), .Y(n3738)
         );
  AND4X1_RVT U3567 ( .A1(n3475), .A2(n3665), .A3(n3743), .A4(n3744), .Y(n3742)
         );
  OR2X1_RVT U3568 ( .A1(n3745), .A2(n3746), .Y(n3665) );
  OR2X1_RVT U3569 ( .A1(n3260), .A2(n3530), .Y(n3475) );
  OR2X1_RVT U3570 ( .A1(n12734), .A2(n12560), .Y(n3530) );
  AND4X1_RVT U3571 ( .A1(n3733), .A2(n3599), .A3(n3722), .A4(n3257), .Y(n3741)
         );
  OR2X1_RVT U3572 ( .A1(n3747), .A2(n3447), .Y(n3257) );
  OR2X1_RVT U3573 ( .A1(n3262), .A2(n3748), .Y(n3722) );
  OR2X1_RVT U3574 ( .A1(n3295), .A2(n254), .Y(n3599) );
  OR2X1_RVT U3575 ( .A1(n3286), .A2(n3749), .Y(n3733) );
  OR2X1_RVT U3576 ( .A1(n12550), .A2(n12570), .Y(n3749) );
  AND4X1_RVT U3577 ( .A1(n3750), .A2(n3751), .A3(n3752), .A4(n3753), .Y(n3740)
         );
  OR2X1_RVT U3578 ( .A1(n3539), .A2(n3754), .Y(n3753) );
  OR2X1_RVT U3579 ( .A1(n12570), .A2(n3319), .Y(n3754) );
  OR2X1_RVT U3580 ( .A1(n3448), .A2(n3755), .Y(n3752) );
  OR2X1_RVT U3581 ( .A1(n12735), .A2(n3336), .Y(n3755) );
  OR2X1_RVT U3582 ( .A1(n3674), .A2(n3756), .Y(n3751) );
  OR2X1_RVT U3583 ( .A1(n3757), .A2(n3333), .Y(n3756) );
  OR2X1_RVT U3584 ( .A1(n12567), .A2(n3758), .Y(n3750) );
  OR2X1_RVT U3585 ( .A1(n3759), .A2(n12550), .Y(n3758) );
  AND2X1_RVT U3586 ( .A1(n3547), .A2(n3760), .Y(n3759) );
  AND2X1_RVT U3587 ( .A1(n3761), .A2(n3762), .Y(n3739) );
  OR2X1_RVT U3588 ( .A1(n3763), .A2(n3314), .Y(n3762) );
  AND2X1_RVT U3589 ( .A1(n3764), .A2(n3765), .Y(n3763) );
  OR2X1_RVT U3590 ( .A1(n12549), .A2(n3507), .Y(n3765) );
  OR2X1_RVT U3591 ( .A1(n12553), .A2(n3582), .Y(n3764) );
  AND2X1_RVT U3592 ( .A1(n3766), .A2(n3767), .Y(n3761) );
  OR2X1_RVT U3593 ( .A1(n3768), .A2(n3353), .Y(n3767) );
  AND2X1_RVT U3594 ( .A1(n3769), .A2(n3770), .Y(n3768) );
  OR2X1_RVT U3595 ( .A1(n12556), .A2(n264), .Y(n3770) );
  NAND2X1_RVT U3596 ( .A1(n3336), .A2(n12727), .Y(n3769) );
  OR2X1_RVT U3597 ( .A1(n3771), .A2(n256), .Y(n3766) );
  AND2X1_RVT U3598 ( .A1(n3560), .A2(n3437), .Y(n3771) );
  OR2X1_RVT U3599 ( .A1(n3286), .A2(n3772), .Y(n3437) );
  OR2X1_RVT U3600 ( .A1(n12738), .A2(n12545), .Y(n3772) );
  AND4X1_RVT U3601 ( .A1(n3454), .A2(n3773), .A3(n3646), .A4(n3774), .Y(n3737)
         );
  AND4X1_RVT U3602 ( .A1(n3775), .A2(n3776), .A3(n3777), .A4(n3778), .Y(n3774)
         );
  OR2X1_RVT U3603 ( .A1(n3417), .A2(n3338), .Y(n3778) );
  OR2X1_RVT U3604 ( .A1(n3355), .A2(n3384), .Y(n3777) );
  OR2X1_RVT U3605 ( .A1(n12726), .A2(n3609), .Y(n3776) );
  OR2X1_RVT U3606 ( .A1(n3333), .A2(n3315), .Y(n3609) );
  OR2X1_RVT U3607 ( .A1(n12734), .A2(n3397), .Y(n3315) );
  OR2X1_RVT U3608 ( .A1(n12559), .A2(n3438), .Y(n3775) );
  OR2X1_RVT U3609 ( .A1(n3319), .A2(n3547), .Y(n3438) );
  OR2X1_RVT U3610 ( .A1(n12543), .A2(n3523), .Y(n3547) );
  AND2X1_RVT U3611 ( .A1(n3779), .A2(n3780), .Y(n3646) );
  OR2X1_RVT U3612 ( .A1(n3781), .A2(n3386), .Y(n3780) );
  OR2X1_RVT U3613 ( .A1(n12569), .A2(n256), .Y(n3781) );
  OR2X1_RVT U3614 ( .A1(n3782), .A2(n3269), .Y(n3779) );
  OR2X1_RVT U3615 ( .A1(n12725), .A2(n3386), .Y(n3269) );
  OR2X1_RVT U3616 ( .A1(n3283), .A2(n3333), .Y(n3782) );
  OR2X1_RVT U3617 ( .A1(n12551), .A2(n3652), .Y(n3773) );
  AND2X1_RVT U3618 ( .A1(n3783), .A2(n3784), .Y(n3454) );
  OR2X1_RVT U3619 ( .A1(n3337), .A2(n3375), .Y(n3784) );
  OR2X1_RVT U3620 ( .A1(n3785), .A2(n3786), .Y(n3783) );
  AND4X1_RVT U3621 ( .A1(n3787), .A2(n3788), .A3(n3789), .A4(n3790), .Y(n3736)
         );
  OR2X1_RVT U3622 ( .A1(n3791), .A2(n3523), .Y(n3790) );
  AND2X1_RVT U3623 ( .A1(n3792), .A2(n3532), .Y(n3791) );
  OR2X1_RVT U3624 ( .A1(n12557), .A2(n3748), .Y(n3532) );
  OR2X1_RVT U3625 ( .A1(n3793), .A2(n12731), .Y(n3789) );
  AND2X1_RVT U3626 ( .A1(n3460), .A2(n3425), .Y(n3793) );
  OR2X1_RVT U3627 ( .A1(n12725), .A2(n3401), .Y(n3425) );
  OR2X1_RVT U3628 ( .A1(n3794), .A2(n3480), .Y(n3788) );
  AND2X1_RVT U3629 ( .A1(n3795), .A2(n3796), .Y(n3794) );
  OR2X1_RVT U3630 ( .A1(n12546), .A2(n3339), .Y(n3796) );
  AND2X1_RVT U3631 ( .A1(n3797), .A2(n3377), .Y(n3795) );
  OR2X1_RVT U3632 ( .A1(n254), .A2(n3336), .Y(n3797) );
  OR2X1_RVT U3633 ( .A1(n3798), .A2(n3277), .Y(n3787) );
  AND2X1_RVT U3634 ( .A1(n3799), .A2(n3800), .Y(n3798) );
  NAND2X1_RVT U3635 ( .A1(n3262), .A2(n3640), .Y(n3800) );
  AND2X1_RVT U3636 ( .A1(n3801), .A2(n3490), .Y(n3799) );
  OR2X1_RVT U3637 ( .A1(n3423), .A2(n3748), .Y(n3490) );
  OR2X1_RVT U3638 ( .A1(n12566), .A2(n3802), .Y(n3801) );
  AND4X1_RVT U3639 ( .A1(n3803), .A2(n3804), .A3(n3805), .A4(n3806), .Y(n3735)
         );
  OR2X1_RVT U3640 ( .A1(n3807), .A2(n3300), .Y(n3806) );
  AND2X1_RVT U3641 ( .A1(n3808), .A2(n3441), .Y(n3807) );
  AND2X1_RVT U3642 ( .A1(n3809), .A2(n3463), .Y(n3808) );
  OR2X1_RVT U3643 ( .A1(n256), .A2(n3786), .Y(n3463) );
  OR2X1_RVT U3644 ( .A1(n12545), .A2(n3397), .Y(n3786) );
  OR2X1_RVT U3645 ( .A1(n3810), .A2(n12562), .Y(n3805) );
  AND2X1_RVT U3646 ( .A1(n3811), .A2(n3812), .Y(n3810) );
  OR2X1_RVT U3647 ( .A1(n3813), .A2(n12723), .Y(n3812) );
  AND2X1_RVT U3648 ( .A1(n3814), .A2(n3815), .Y(n3813) );
  OR2X1_RVT U3649 ( .A1(n12544), .A2(n3674), .Y(n3815) );
  OR2X1_RVT U3650 ( .A1(n12730), .A2(n3320), .Y(n3814) );
  AND2X1_RVT U3651 ( .A1(n3816), .A2(n3817), .Y(n3811) );
  OR2X1_RVT U3652 ( .A1(n3286), .A2(n3818), .Y(n3816) );
  OR2X1_RVT U3653 ( .A1(n3819), .A2(n3320), .Y(n3804) );
  AND4X1_RVT U3654 ( .A1(n3820), .A2(n3821), .A3(n3822), .A4(n3286), .Y(n3819)
         );
  OR2X1_RVT U3655 ( .A1(n12731), .A2(n3336), .Y(n3822) );
  OR2X1_RVT U3656 ( .A1(n12556), .A2(n3355), .Y(n3821) );
  OR2X1_RVT U3657 ( .A1(n3408), .A2(n3386), .Y(n3820) );
  OR2X1_RVT U3658 ( .A1(n3823), .A2(n3262), .Y(n3803) );
  AND4X1_RVT U3659 ( .A1(n3687), .A2(n3824), .A3(n3485), .A4(n3401), .Y(n3823)
         );
  OR2X1_RVT U3660 ( .A1(n3355), .A2(n3818), .Y(n3485) );
  OR2X1_RVT U3661 ( .A1(n3523), .A2(n3730), .Y(n3824) );
  OR2X1_RVT U3662 ( .A1(n12550), .A2(n3488), .Y(n3687) );
  AND4X1_RVT U3663 ( .A1(n3826), .A2(n3827), .A3(n3828), .A4(n3829), .Y(n3825)
         );
  AND4X1_RVT U3664 ( .A1(n3338), .A2(n3574), .A3(n3830), .A4(n3831), .Y(n3829)
         );
  AND4X1_RVT U3665 ( .A1(n3653), .A2(n3598), .A3(n3743), .A4(n3744), .Y(n3831)
         );
  OR2X1_RVT U3666 ( .A1(n3746), .A2(n3259), .Y(n3744) );
  OR2X1_RVT U3667 ( .A1(n12729), .A2(n3377), .Y(n3259) );
  OR2X1_RVT U3668 ( .A1(n3276), .A2(n3785), .Y(n3743) );
  OR2X1_RVT U3669 ( .A1(n12734), .A2(n12564), .Y(n3785) );
  OR2X1_RVT U3670 ( .A1(n12723), .A2(n3397), .Y(n3276) );
  OR2X1_RVT U3671 ( .A1(n12735), .A2(n3295), .Y(n3598) );
  OR2X1_RVT U3672 ( .A1(n12573), .A2(n12557), .Y(n3295) );
  OR2X1_RVT U3673 ( .A1(n3417), .A2(n3832), .Y(n3653) );
  OR2X1_RVT U3674 ( .A1(n12564), .A2(n3321), .Y(n3832) );
  OR2X1_RVT U3675 ( .A1(n3319), .A2(n3833), .Y(n3830) );
  OR2X1_RVT U3676 ( .A1(n3447), .A2(n12555), .Y(n3833) );
  OR2X1_RVT U3677 ( .A1(n3386), .A2(n3834), .Y(n3574) );
  OR2X1_RVT U3678 ( .A1(n3320), .A2(n12562), .Y(n3834) );
  OR2X1_RVT U3679 ( .A1(n12727), .A2(n3745), .Y(n3338) );
  OR2X1_RVT U3680 ( .A1(n12557), .A2(n3337), .Y(n3745) );
  AND4X1_RVT U3681 ( .A1(n3835), .A2(n3836), .A3(n3837), .A4(n3838), .Y(n3828)
         );
  AND4X1_RVT U3682 ( .A1(n3839), .A2(n3840), .A3(n3841), .A4(n3842), .Y(n3838)
         );
  OR2X1_RVT U3683 ( .A1(n3353), .A2(n3843), .Y(n3842) );
  OR2X1_RVT U3684 ( .A1(n12546), .A2(n3423), .Y(n3843) );
  OR2X1_RVT U3685 ( .A1(n3336), .A2(n3844), .Y(n3841) );
  OR2X1_RVT U3686 ( .A1(n3845), .A2(n3300), .Y(n3844) );
  AND2X1_RVT U3687 ( .A1(n3279), .A2(n3339), .Y(n3845) );
  OR2X1_RVT U3688 ( .A1(n3846), .A2(n3847), .Y(n3840) );
  AND2X1_RVT U3689 ( .A1(n3494), .A2(n3450), .Y(n3846) );
  OR2X1_RVT U3690 ( .A1(n12728), .A2(n264), .Y(n3450) );
  OR2X1_RVT U3691 ( .A1(n12724), .A2(n12567), .Y(n3494) );
  OR2X1_RVT U3692 ( .A1(n3848), .A2(n3334), .Y(n3839) );
  AND2X1_RVT U3693 ( .A1(n3730), .A2(n3849), .Y(n3848) );
  OR2X1_RVT U3694 ( .A1(n12726), .A2(n256), .Y(n3849) );
  OR2X1_RVT U3695 ( .A1(n3850), .A2(n12569), .Y(n3837) );
  AND2X1_RVT U3696 ( .A1(n3721), .A2(n3851), .Y(n3850) );
  OR2X1_RVT U3697 ( .A1(n3327), .A2(n3674), .Y(n3851) );
  OR2X1_RVT U3698 ( .A1(n12550), .A2(n3539), .Y(n3721) );
  OR2X1_RVT U3699 ( .A1(n12730), .A2(n3327), .Y(n3539) );
  OR2X1_RVT U3700 ( .A1(n3852), .A2(n3488), .Y(n3836) );
  AND2X1_RVT U3701 ( .A1(n3441), .A2(n3713), .Y(n3852) );
  OR2X1_RVT U3702 ( .A1(n3297), .A2(n3386), .Y(n3441) );
  OR2X1_RVT U3703 ( .A1(n3853), .A2(n3377), .Y(n3835) );
  AND2X1_RVT U3704 ( .A1(n3340), .A2(n3342), .Y(n3853) );
  AND4X1_RVT U3705 ( .A1(n3854), .A2(n3855), .A3(n3856), .A4(n3857), .Y(n3827)
         );
  AND4X1_RVT U3706 ( .A1(n3858), .A2(n3859), .A3(n3860), .A4(n3861), .Y(n3857)
         );
  OR2X1_RVT U3707 ( .A1(n3862), .A2(n12553), .Y(n3861) );
  AND2X1_RVT U3708 ( .A1(n3268), .A2(n3560), .Y(n3862) );
  OR2X1_RVT U3709 ( .A1(n3417), .A2(n3448), .Y(n3560) );
  OR2X1_RVT U3710 ( .A1(n12556), .A2(n3300), .Y(n3448) );
  OR2X1_RVT U3711 ( .A1(n12560), .A2(n3863), .Y(n3268) );
  OR2X1_RVT U3712 ( .A1(n12543), .A2(n12549), .Y(n3863) );
  OR2X1_RVT U3713 ( .A1(n3864), .A2(n12567), .Y(n3860) );
  AND2X1_RVT U3714 ( .A1(n3577), .A2(n3865), .Y(n3864) );
  OR2X1_RVT U3715 ( .A1(n12572), .A2(n254), .Y(n3865) );
  OR2X1_RVT U3716 ( .A1(n12570), .A2(n3384), .Y(n3577) );
  OR2X1_RVT U3717 ( .A1(n3866), .A2(n12548), .Y(n3859) );
  AND2X1_RVT U3718 ( .A1(n3595), .A2(n3867), .Y(n3866) );
  OR2X1_RVT U3719 ( .A1(n12573), .A2(n3320), .Y(n3867) );
  OR2X1_RVT U3720 ( .A1(n3262), .A2(n3868), .Y(n3595) );
  OR2X1_RVT U3721 ( .A1(n3869), .A2(n3321), .Y(n3858) );
  AND2X1_RVT U3722 ( .A1(n3870), .A2(n3871), .Y(n3869) );
  OR2X1_RVT U3723 ( .A1(n3377), .A2(n12570), .Y(n3871) );
  AND2X1_RVT U3724 ( .A1(n3872), .A2(n3353), .Y(n3870) );
  OR2X1_RVT U3725 ( .A1(n3339), .A2(n3300), .Y(n3353) );
  OR2X1_RVT U3726 ( .A1(n12545), .A2(n3384), .Y(n3872) );
  OR2X1_RVT U3727 ( .A1(n12738), .A2(n3339), .Y(n3384) );
  OR2X1_RVT U3728 ( .A1(n3873), .A2(n3397), .Y(n3856) );
  AND4X1_RVT U3729 ( .A1(n3874), .A2(n3875), .A3(n3550), .A4(n3460), .Y(n3873)
         );
  OR2X1_RVT U3730 ( .A1(n3523), .A2(n3623), .Y(n3460) );
  OR2X1_RVT U3731 ( .A1(n3355), .A2(n3802), .Y(n3550) );
  OR2X1_RVT U3732 ( .A1(n12551), .A2(n12544), .Y(n3802) );
  OR2X1_RVT U3733 ( .A1(n256), .A2(n3277), .Y(n3875) );
  OR2X1_RVT U3734 ( .A1(n254), .A2(n12570), .Y(n3874) );
  OR2X1_RVT U3735 ( .A1(n3876), .A2(n3333), .Y(n3855) );
  AND2X1_RVT U3736 ( .A1(n3877), .A2(n3354), .Y(n3876) );
  AND2X1_RVT U3737 ( .A1(n3809), .A2(n3604), .Y(n3877) );
  OR2X1_RVT U3738 ( .A1(n3878), .A2(n12735), .Y(n3604) );
  AND2X1_RVT U3739 ( .A1(n3375), .A2(n3879), .Y(n3878) );
  OR2X1_RVT U3740 ( .A1(n12548), .A2(n3262), .Y(n3879) );
  OR2X1_RVT U3741 ( .A1(n3423), .A2(n3561), .Y(n3809) );
  OR2X1_RVT U3742 ( .A1(n3408), .A2(n3297), .Y(n3561) );
  OR2X1_RVT U3743 ( .A1(n3880), .A2(n3401), .Y(n3854) );
  AND2X1_RVT U3744 ( .A1(n3881), .A2(n12556), .Y(n3880) );
  AND2X1_RVT U3745 ( .A1(n3882), .A2(n3582), .Y(n3881) );
  OR2X1_RVT U3746 ( .A1(n3423), .A2(n3523), .Y(n3882) );
  AND4X1_RVT U3747 ( .A1(n3883), .A2(n3884), .A3(n3885), .A4(n3886), .Y(n3826)
         );
  AND2X1_RVT U3748 ( .A1(n3887), .A2(n3888), .Y(n3886) );
  OR2X1_RVT U3749 ( .A1(n12731), .A2(n3503), .Y(n3888) );
  OR2X1_RVT U3750 ( .A1(n12564), .A2(n3889), .Y(n3503) );
  OR2X1_RVT U3751 ( .A1(n3319), .A2(n3408), .Y(n3889) );
  AND2X1_RVT U3752 ( .A1(n3890), .A2(n3891), .Y(n3887) );
  OR2X1_RVT U3753 ( .A1(n3292), .A2(n3303), .Y(n3891) );
  OR2X1_RVT U3754 ( .A1(n3336), .A2(n3531), .Y(n3303) );
  OR2X1_RVT U3755 ( .A1(n12727), .A2(n3297), .Y(n3531) );
  OR2X1_RVT U3756 ( .A1(n3339), .A2(n3416), .Y(n3890) );
  OR2X1_RVT U3757 ( .A1(n3327), .A2(n3892), .Y(n3416) );
  OR2X1_RVT U3758 ( .A1(n3327), .A2(n3507), .Y(n3885) );
  OR2X1_RVT U3759 ( .A1(n256), .A2(n12566), .Y(n3507) );
  OR2X1_RVT U3760 ( .A1(n3893), .A2(n3283), .Y(n3884) );
  AND4X1_RVT U3761 ( .A1(n3894), .A2(n3895), .A3(n3896), .A4(n3897), .Y(n3893)
         );
  OR2X1_RVT U3762 ( .A1(n12725), .A2(n3898), .Y(n3896) );
  OR2X1_RVT U3763 ( .A1(n3899), .A2(n12732), .Y(n3898) );
  AND2X1_RVT U3764 ( .A1(n3334), .A2(n3900), .Y(n3899) );
  OR2X1_RVT U3765 ( .A1(n12559), .A2(n3901), .Y(n3895) );
  OR2X1_RVT U3766 ( .A1(n3640), .A2(n3277), .Y(n3901) );
  OR2X1_RVT U3767 ( .A1(n3260), .A2(n3286), .Y(n3894) );
  OR2X1_RVT U3768 ( .A1(n12729), .A2(n3386), .Y(n3286) );
  OR2X1_RVT U3769 ( .A1(n3760), .A2(n3674), .Y(n3883) );
  OR2X1_RVT U3770 ( .A1(n12575), .A2(n3297), .Y(n3674) );
  AND4X1_RVT U3771 ( .A1(n3903), .A2(n3904), .A3(n3905), .A4(n3906), .Y(n3902)
         );
  AND4X1_RVT U3772 ( .A1(n2758), .A2(n2994), .A3(n3907), .A4(n3908), .Y(n3906)
         );
  AND4X1_RVT U3773 ( .A1(n3073), .A2(n3018), .A3(n3163), .A4(n3164), .Y(n3908)
         );
  OR2X1_RVT U3774 ( .A1(n3166), .A2(n2679), .Y(n3164) );
  OR2X1_RVT U3775 ( .A1(n12884), .A2(n2797), .Y(n2679) );
  OR2X1_RVT U3776 ( .A1(n2696), .A2(n3205), .Y(n3163) );
  OR2X1_RVT U3777 ( .A1(n12889), .A2(n12498), .Y(n3205) );
  OR2X1_RVT U3778 ( .A1(n12878), .A2(n2817), .Y(n2696) );
  OR2X1_RVT U3779 ( .A1(n12890), .A2(n2715), .Y(n3018) );
  OR2X1_RVT U3780 ( .A1(n12507), .A2(n12491), .Y(n2715) );
  OR2X1_RVT U3781 ( .A1(n2837), .A2(n3909), .Y(n3073) );
  OR2X1_RVT U3782 ( .A1(n12498), .A2(n2741), .Y(n3909) );
  OR2X1_RVT U3783 ( .A1(n2739), .A2(n3910), .Y(n3907) );
  OR2X1_RVT U3784 ( .A1(n2867), .A2(n12489), .Y(n3910) );
  OR2X1_RVT U3785 ( .A1(n2806), .A2(n3911), .Y(n2994) );
  OR2X1_RVT U3786 ( .A1(n2740), .A2(n12496), .Y(n3911) );
  OR2X1_RVT U3787 ( .A1(n12882), .A2(n3165), .Y(n2758) );
  OR2X1_RVT U3788 ( .A1(n12491), .A2(n2757), .Y(n3165) );
  AND4X1_RVT U3789 ( .A1(n3912), .A2(n3913), .A3(n3914), .A4(n3915), .Y(n3905)
         );
  AND4X1_RVT U3790 ( .A1(n3916), .A2(n3917), .A3(n3918), .A4(n3919), .Y(n3915)
         );
  OR2X1_RVT U3791 ( .A1(n2773), .A2(n3920), .Y(n3919) );
  OR2X1_RVT U3792 ( .A1(n12480), .A2(n2843), .Y(n3920) );
  OR2X1_RVT U3793 ( .A1(n2756), .A2(n3921), .Y(n3918) );
  OR2X1_RVT U3794 ( .A1(n3922), .A2(n2720), .Y(n3921) );
  AND2X1_RVT U3795 ( .A1(n2699), .A2(n2759), .Y(n3922) );
  OR2X1_RVT U3796 ( .A1(n3923), .A2(n3924), .Y(n3917) );
  AND2X1_RVT U3797 ( .A1(n2914), .A2(n2870), .Y(n3923) );
  OR2X1_RVT U3798 ( .A1(n12883), .A2(n59), .Y(n2870) );
  OR2X1_RVT U3799 ( .A1(n12879), .A2(n12501), .Y(n2914) );
  OR2X1_RVT U3800 ( .A1(n3925), .A2(n2754), .Y(n3916) );
  AND2X1_RVT U3801 ( .A1(n3150), .A2(n3926), .Y(n3925) );
  OR2X1_RVT U3802 ( .A1(n12881), .A2(n51), .Y(n3926) );
  OR2X1_RVT U3803 ( .A1(n3927), .A2(n12503), .Y(n3914) );
  AND2X1_RVT U3804 ( .A1(n3141), .A2(n3928), .Y(n3927) );
  OR2X1_RVT U3805 ( .A1(n2747), .A2(n3094), .Y(n3928) );
  OR2X1_RVT U3806 ( .A1(n12484), .A2(n2959), .Y(n3141) );
  OR2X1_RVT U3807 ( .A1(n12885), .A2(n2747), .Y(n2959) );
  OR2X1_RVT U3808 ( .A1(n3929), .A2(n2908), .Y(n3913) );
  AND2X1_RVT U3809 ( .A1(n2861), .A2(n3133), .Y(n3929) );
  OR2X1_RVT U3810 ( .A1(n2717), .A2(n2806), .Y(n2861) );
  OR2X1_RVT U3811 ( .A1(n3930), .A2(n2797), .Y(n3912) );
  AND2X1_RVT U3812 ( .A1(n2760), .A2(n2762), .Y(n3930) );
  AND4X1_RVT U3813 ( .A1(n3931), .A2(n3932), .A3(n3933), .A4(n3934), .Y(n3904)
         );
  AND4X1_RVT U3814 ( .A1(n3935), .A2(n3936), .A3(n3937), .A4(n3938), .Y(n3934)
         );
  OR2X1_RVT U3815 ( .A1(n3939), .A2(n12487), .Y(n3938) );
  AND2X1_RVT U3816 ( .A1(n2688), .A2(n2980), .Y(n3939) );
  OR2X1_RVT U3817 ( .A1(n2837), .A2(n2868), .Y(n2980) );
  OR2X1_RVT U3818 ( .A1(n12490), .A2(n2720), .Y(n2868) );
  OR2X1_RVT U3819 ( .A1(n12494), .A2(n3940), .Y(n2688) );
  OR2X1_RVT U3820 ( .A1(n12477), .A2(n12483), .Y(n3940) );
  OR2X1_RVT U3821 ( .A1(n3941), .A2(n12501), .Y(n3937) );
  AND2X1_RVT U3822 ( .A1(n2997), .A2(n3942), .Y(n3941) );
  OR2X1_RVT U3823 ( .A1(n12506), .A2(n49), .Y(n3942) );
  OR2X1_RVT U3824 ( .A1(n12504), .A2(n2804), .Y(n2997) );
  OR2X1_RVT U3825 ( .A1(n3943), .A2(n12482), .Y(n3936) );
  AND2X1_RVT U3826 ( .A1(n3015), .A2(n3944), .Y(n3943) );
  OR2X1_RVT U3827 ( .A1(n12507), .A2(n2740), .Y(n3944) );
  OR2X1_RVT U3828 ( .A1(n2682), .A2(n3945), .Y(n3015) );
  OR2X1_RVT U3829 ( .A1(n3946), .A2(n2741), .Y(n3935) );
  AND2X1_RVT U3830 ( .A1(n3947), .A2(n3948), .Y(n3946) );
  OR2X1_RVT U3831 ( .A1(n2797), .A2(n12504), .Y(n3948) );
  AND2X1_RVT U3832 ( .A1(n3949), .A2(n2773), .Y(n3947) );
  OR2X1_RVT U3833 ( .A1(n2759), .A2(n2720), .Y(n2773) );
  OR2X1_RVT U3834 ( .A1(n12479), .A2(n2804), .Y(n3949) );
  OR2X1_RVT U3835 ( .A1(n12893), .A2(n2759), .Y(n2804) );
  OR2X1_RVT U3836 ( .A1(n3950), .A2(n2817), .Y(n3933) );
  AND4X1_RVT U3837 ( .A1(n3951), .A2(n3952), .A3(n2970), .A4(n2880), .Y(n3950)
         );
  OR2X1_RVT U3838 ( .A1(n2943), .A2(n3043), .Y(n2880) );
  OR2X1_RVT U3839 ( .A1(n2775), .A2(n3222), .Y(n2970) );
  OR2X1_RVT U3840 ( .A1(n12485), .A2(n12478), .Y(n3222) );
  OR2X1_RVT U3841 ( .A1(n51), .A2(n2697), .Y(n3952) );
  OR2X1_RVT U3842 ( .A1(n49), .A2(n12504), .Y(n3951) );
  OR2X1_RVT U3843 ( .A1(n3953), .A2(n2753), .Y(n3932) );
  AND2X1_RVT U3844 ( .A1(n3954), .A2(n2774), .Y(n3953) );
  AND2X1_RVT U3845 ( .A1(n3229), .A2(n3024), .Y(n3954) );
  OR2X1_RVT U3846 ( .A1(n3955), .A2(n12890), .Y(n3024) );
  AND2X1_RVT U3847 ( .A1(n2795), .A2(n3956), .Y(n3955) );
  OR2X1_RVT U3848 ( .A1(n12482), .A2(n2682), .Y(n3956) );
  OR2X1_RVT U3849 ( .A1(n2843), .A2(n2981), .Y(n3229) );
  OR2X1_RVT U3850 ( .A1(n2828), .A2(n2717), .Y(n2981) );
  OR2X1_RVT U3851 ( .A1(n3957), .A2(n2821), .Y(n3931) );
  AND2X1_RVT U3852 ( .A1(n3958), .A2(n12490), .Y(n3957) );
  AND2X1_RVT U3853 ( .A1(n3959), .A2(n3002), .Y(n3958) );
  OR2X1_RVT U3854 ( .A1(n2843), .A2(n2943), .Y(n3959) );
  AND4X1_RVT U3855 ( .A1(n3960), .A2(n3961), .A3(n3962), .A4(n3963), .Y(n3903)
         );
  AND2X1_RVT U3856 ( .A1(n3964), .A2(n3965), .Y(n3963) );
  OR2X1_RVT U3857 ( .A1(n12886), .A2(n2923), .Y(n3965) );
  OR2X1_RVT U3858 ( .A1(n12498), .A2(n3966), .Y(n2923) );
  OR2X1_RVT U3859 ( .A1(n2739), .A2(n2828), .Y(n3966) );
  AND2X1_RVT U3860 ( .A1(n3967), .A2(n3968), .Y(n3964) );
  OR2X1_RVT U3861 ( .A1(n2712), .A2(n2723), .Y(n3968) );
  OR2X1_RVT U3862 ( .A1(n2756), .A2(n2951), .Y(n2723) );
  OR2X1_RVT U3863 ( .A1(n12882), .A2(n2717), .Y(n2951) );
  OR2X1_RVT U3864 ( .A1(n2759), .A2(n2836), .Y(n3967) );
  OR2X1_RVT U3865 ( .A1(n2747), .A2(n3969), .Y(n2836) );
  OR2X1_RVT U3866 ( .A1(n2747), .A2(n2927), .Y(n3962) );
  OR2X1_RVT U3867 ( .A1(n51), .A2(n12500), .Y(n2927) );
  OR2X1_RVT U3868 ( .A1(n3970), .A2(n2703), .Y(n3961) );
  AND4X1_RVT U3869 ( .A1(n3971), .A2(n3972), .A3(n3973), .A4(n3974), .Y(n3970)
         );
  OR2X1_RVT U3870 ( .A1(n12880), .A2(n3975), .Y(n3973) );
  OR2X1_RVT U3871 ( .A1(n3976), .A2(n12887), .Y(n3975) );
  AND2X1_RVT U3872 ( .A1(n2754), .A2(n3977), .Y(n3976) );
  OR2X1_RVT U3873 ( .A1(n12493), .A2(n3978), .Y(n3972) );
  OR2X1_RVT U3874 ( .A1(n3060), .A2(n2697), .Y(n3978) );
  OR2X1_RVT U3875 ( .A1(n2680), .A2(n2706), .Y(n3971) );
  OR2X1_RVT U3876 ( .A1(n12884), .A2(n2806), .Y(n2706) );
  OR2X1_RVT U3877 ( .A1(n3180), .A2(n3094), .Y(n3960) );
  OR2X1_RVT U3878 ( .A1(n12509), .A2(n2717), .Y(n3094) );
  AND4X1_RVT U3879 ( .A1(n3980), .A2(n3981), .A3(n3982), .A4(n3983), .Y(n3979)
         );
  AND4X1_RVT U3880 ( .A1(n3984), .A2(n3985), .A3(n3986), .A4(n3987), .Y(n3983)
         );
  AND4X1_RVT U3881 ( .A1(n3988), .A2(n3989), .A3(n3990), .A4(n3991), .Y(n3987)
         );
  OR2X1_RVT U3882 ( .A1(n3748), .A2(n3892), .Y(n3991) );
  OR2X1_RVT U3883 ( .A1(n12728), .A2(n12569), .Y(n3892) );
  OR2X1_RVT U3884 ( .A1(n12543), .A2(n12553), .Y(n3748) );
  OR2X1_RVT U3885 ( .A1(n3992), .A2(n3334), .Y(n3990) );
  AND2X1_RVT U3886 ( .A1(n3280), .A2(n3847), .Y(n3992) );
  OR2X1_RVT U3887 ( .A1(n256), .A2(n3993), .Y(n3280) );
  OR2X1_RVT U3888 ( .A1(n12543), .A2(n12725), .Y(n3993) );
  OR2X1_RVT U3889 ( .A1(n3994), .A2(n3262), .Y(n3989) );
  OR2X1_RVT U3890 ( .A1(n12557), .A2(n3423), .Y(n3262) );
  AND2X1_RVT U3891 ( .A1(n3398), .A2(n3995), .Y(n3994) );
  OR2X1_RVT U3892 ( .A1(n3277), .A2(n3479), .Y(n3995) );
  OR2X1_RVT U3893 ( .A1(n12561), .A2(n12549), .Y(n3277) );
  OR2X1_RVT U3894 ( .A1(n3523), .A2(n3996), .Y(n3398) );
  OR2X1_RVT U3895 ( .A1(n12736), .A2(n12564), .Y(n3996) );
  OR2X1_RVT U3896 ( .A1(n3997), .A2(n3321), .Y(n3988) );
  AND2X1_RVT U3897 ( .A1(n3718), .A2(n3998), .Y(n3997) );
  OR2X1_RVT U3898 ( .A1(n3999), .A2(n12725), .Y(n3998) );
  AND2X1_RVT U3899 ( .A1(n3377), .A2(n3730), .Y(n3999) );
  OR2X1_RVT U3900 ( .A1(n12733), .A2(n3339), .Y(n3730) );
  OR2X1_RVT U3901 ( .A1(n12570), .A2(n4000), .Y(n3718) );
  OR2X1_RVT U3902 ( .A1(n12738), .A2(n12734), .Y(n4000) );
  OR2X1_RVT U3903 ( .A1(n4001), .A2(n12548), .Y(n3986) );
  AND2X1_RVT U3904 ( .A1(n4002), .A2(n4003), .Y(n4001) );
  OR2X1_RVT U3905 ( .A1(n4004), .A2(n3423), .Y(n4003) );
  AND2X1_RVT U3906 ( .A1(n3488), .A2(n4005), .Y(n4004) );
  OR2X1_RVT U3907 ( .A1(n3279), .A2(n3401), .Y(n4002) );
  OR2X1_RVT U3908 ( .A1(n12562), .A2(n3337), .Y(n3401) );
  OR2X1_RVT U3909 ( .A1(n4006), .A2(n12734), .Y(n3985) );
  AND2X1_RVT U3910 ( .A1(n3493), .A2(n3652), .Y(n4006) );
  OR2X1_RVT U3911 ( .A1(n12560), .A2(n4007), .Y(n3652) );
  OR2X1_RVT U3912 ( .A1(n3333), .A2(n12549), .Y(n4007) );
  OR2X1_RVT U3913 ( .A1(n3279), .A2(n3760), .Y(n3493) );
  OR2X1_RVT U3914 ( .A1(n12549), .A2(n12564), .Y(n3760) );
  OR2X1_RVT U3915 ( .A1(n4008), .A2(n12546), .Y(n3984) );
  AND2X1_RVT U3916 ( .A1(n3533), .A2(n4009), .Y(n4008) );
  OR2X1_RVT U3917 ( .A1(n3747), .A2(n3327), .Y(n4009) );
  OR2X1_RVT U3918 ( .A1(n3386), .A2(n3868), .Y(n3533) );
  OR2X1_RVT U3919 ( .A1(n12733), .A2(n256), .Y(n3868) );
  AND2X1_RVT U3920 ( .A1(n12550), .A2(n12736), .Y(n3629) );
  AND4X1_RVT U3921 ( .A1(n4010), .A2(n4011), .A3(n4012), .A4(n4013), .Y(n3982)
         );
  AND4X1_RVT U3922 ( .A1(n4014), .A2(n4015), .A3(n4016), .A4(n4017), .Y(n4013)
         );
  OR2X1_RVT U3923 ( .A1(n4018), .A2(n12555), .Y(n4017) );
  AND2X1_RVT U3924 ( .A1(n3520), .A2(n3591), .Y(n4018) );
  OR2X1_RVT U3925 ( .A1(n3336), .A2(n3847), .Y(n3591) );
  OR2X1_RVT U3926 ( .A1(n12736), .A2(n3333), .Y(n3847) );
  OR2X1_RVT U3927 ( .A1(n12723), .A2(n12545), .Y(n3336) );
  OR2X1_RVT U3928 ( .A1(n12546), .A2(n3623), .Y(n3520) );
  OR2X1_RVT U3929 ( .A1(n12550), .A2(n12564), .Y(n3623) );
  OR2X1_RVT U3930 ( .A1(n4019), .A2(n12732), .Y(n4016) );
  AND2X1_RVT U3931 ( .A1(n3682), .A2(n4020), .Y(n4019) );
  OR2X1_RVT U3932 ( .A1(n3640), .A2(n3350), .Y(n4020) );
  OR2X1_RVT U3933 ( .A1(n3523), .A2(n4021), .Y(n3350) );
  OR2X1_RVT U3934 ( .A1(n12575), .A2(n12551), .Y(n4021) );
  OR2X1_RVT U3935 ( .A1(n12559), .A2(n4022), .Y(n3682) );
  OR2X1_RVT U3936 ( .A1(n3523), .A2(n3319), .Y(n4022) );
  OR2X1_RVT U3937 ( .A1(n4023), .A2(n12738), .Y(n4015) );
  AND2X1_RVT U3938 ( .A1(n3628), .A2(n3557), .Y(n4023) );
  OR2X1_RVT U3939 ( .A1(n3339), .A2(n3375), .Y(n3557) );
  OR2X1_RVT U3940 ( .A1(n12730), .A2(n3523), .Y(n3375) );
  OR2X1_RVT U3941 ( .A1(n3747), .A2(n3355), .Y(n3628) );
  OR2X1_RVT U3942 ( .A1(n12556), .A2(n12735), .Y(n3747) );
  OR2X1_RVT U3943 ( .A1(n4024), .A2(n3397), .Y(n4014) );
  AND2X1_RVT U3944 ( .A1(n4025), .A2(n4026), .Y(n4024) );
  OR2X1_RVT U3945 ( .A1(n3319), .A2(n3746), .Y(n4026) );
  OR2X1_RVT U3946 ( .A1(n12732), .A2(n264), .Y(n3746) );
  AND2X1_RVT U3947 ( .A1(n4027), .A2(n3614), .Y(n4025) );
  OR2X1_RVT U3948 ( .A1(n3327), .A2(n4028), .Y(n3614) );
  OR2X1_RVT U3949 ( .A1(n12572), .A2(n12551), .Y(n4028) );
  OR2X1_RVT U3950 ( .A1(n3383), .A2(n3320), .Y(n4012) );
  OR2X1_RVT U3951 ( .A1(n12725), .A2(n3279), .Y(n3383) );
  OR2X1_RVT U3952 ( .A1(n4029), .A2(n3283), .Y(n4011) );
  AND2X1_RVT U3953 ( .A1(n4030), .A2(n3464), .Y(n4029) );
  AND2X1_RVT U3954 ( .A1(n4031), .A2(n4032), .Y(n3464) );
  OR2X1_RVT U3955 ( .A1(n12560), .A2(n3488), .Y(n4032) );
  OR2X1_RVT U3956 ( .A1(n3386), .A2(n3260), .Y(n4031) );
  OR2X1_RVT U3957 ( .A1(n12545), .A2(n3333), .Y(n3260) );
  AND2X1_RVT U3958 ( .A1(n4033), .A2(n3650), .Y(n4030) );
  OR2X1_RVT U3959 ( .A1(n3417), .A2(n3900), .Y(n3650) );
  OR2X1_RVT U3960 ( .A1(n12727), .A2(n254), .Y(n3900) );
  OR2X1_RVT U3961 ( .A1(n3279), .A2(n3446), .Y(n4033) );
  OR2X1_RVT U3962 ( .A1(n12544), .A2(n4034), .Y(n3446) );
  OR2X1_RVT U3963 ( .A1(n12723), .A2(n12573), .Y(n4034) );
  OR2X1_RVT U3964 ( .A1(n4035), .A2(n12723), .Y(n4010) );
  AND4X1_RVT U3965 ( .A1(n4036), .A2(n4037), .A3(n4038), .A4(n3792), .Y(n4035)
         );
  OR2X1_RVT U3966 ( .A1(n3333), .A2(n3713), .Y(n3792) );
  OR2X1_RVT U3967 ( .A1(n12728), .A2(n12734), .Y(n3713) );
  OR2X1_RVT U3968 ( .A1(n3333), .A2(n4039), .Y(n4038) );
  OR2X1_RVT U3969 ( .A1(n12550), .A2(n12555), .Y(n4039) );
  OR2X1_RVT U3970 ( .A1(n12733), .A2(n3292), .Y(n3333) );
  OR2X1_RVT U3971 ( .A1(n4040), .A2(n3414), .Y(n4037) );
  OR2X1_RVT U3972 ( .A1(n12544), .A2(n3258), .Y(n3414) );
  AND2X1_RVT U3973 ( .A1(n3397), .A2(n4041), .Y(n4040) );
  OR2X1_RVT U3974 ( .A1(n12731), .A2(n3297), .Y(n4041) );
  OR2X1_RVT U3975 ( .A1(n12727), .A2(n12555), .Y(n3397) );
  OR2X1_RVT U3976 ( .A1(n12729), .A2(n4005), .Y(n4036) );
  OR2X1_RVT U3977 ( .A1(n12733), .A2(n3337), .Y(n4005) );
  OR2X1_RVT U3978 ( .A1(n3283), .A2(n254), .Y(n3337) );
  AND4X1_RVT U3979 ( .A1(n4042), .A2(n4043), .A3(n4044), .A4(n4045), .Y(n3981)
         );
  AND4X1_RVT U3980 ( .A1(n4046), .A2(n4047), .A3(n4048), .A4(n4049), .Y(n4045)
         );
  OR2X1_RVT U3981 ( .A1(n3355), .A2(n3482), .Y(n4049) );
  OR2X1_RVT U3982 ( .A1(n12557), .A2(n3377), .Y(n3482) );
  OR2X1_RVT U3983 ( .A1(n12561), .A2(n3523), .Y(n3355) );
  OR2X1_RVT U3984 ( .A1(n3342), .A2(n3818), .Y(n4048) );
  OR2X1_RVT U3985 ( .A1(n12737), .A2(n12544), .Y(n3818) );
  OR2X1_RVT U3986 ( .A1(n3408), .A2(n3334), .Y(n3342) );
  OR2X1_RVT U3987 ( .A1(n3327), .A2(n3354), .Y(n4047) );
  OR2X1_RVT U3988 ( .A1(n12553), .A2(n12566), .Y(n3354) );
  OR2X1_RVT U3989 ( .A1(n12543), .A2(n12724), .Y(n3327) );
  OR2X1_RVT U3990 ( .A1(n264), .A2(n3693), .Y(n4046) );
  OR2X1_RVT U3991 ( .A1(n12551), .A2(n3480), .Y(n3693) );
  OR2X1_RVT U3992 ( .A1(n3297), .A2(n3727), .Y(n4044) );
  OR2X1_RVT U3993 ( .A1(n264), .A2(n4050), .Y(n3727) );
  OR2X1_RVT U3994 ( .A1(n12730), .A2(n12564), .Y(n4050) );
  AND2X1_RVT U3995 ( .A1(n12545), .A2(n12548), .Y(n3757) );
  OR2X1_RVT U3996 ( .A1(n3339), .A2(n3287), .Y(n4043) );
  OR2X1_RVT U3997 ( .A1(n12573), .A2(n4051), .Y(n3287) );
  OR2X1_RVT U3998 ( .A1(n12731), .A2(n12723), .Y(n4051) );
  OR2X1_RVT U3999 ( .A1(n12550), .A2(n3319), .Y(n3339) );
  OR2X1_RVT U4000 ( .A1(n3386), .A2(n4027), .Y(n4042) );
  OR2X1_RVT U4001 ( .A1(n12546), .A2(n3341), .Y(n4027) );
  OR2X1_RVT U4002 ( .A1(n12733), .A2(n12734), .Y(n3341) );
  AND4X1_RVT U4003 ( .A1(n4052), .A2(n3452), .A3(n4053), .A4(n4054), .Y(n3980)
         );
  OR2X1_RVT U4004 ( .A1(n12550), .A2(n3897), .Y(n4054) );
  OR2X1_RVT U4005 ( .A1(n12729), .A2(n3447), .Y(n3897) );
  OR2X1_RVT U4006 ( .A1(n12548), .A2(n3488), .Y(n3447) );
  OR2X1_RVT U4007 ( .A1(n12543), .A2(n3314), .Y(n3488) );
  AND2X1_RVT U4008 ( .A1(n4055), .A2(n4056), .Y(n4053) );
  OR2X1_RVT U4009 ( .A1(n12572), .A2(n3817), .Y(n4056) );
  OR2X1_RVT U4010 ( .A1(n3386), .A2(n3479), .Y(n3817) );
  OR2X1_RVT U4011 ( .A1(n12550), .A2(n12544), .Y(n3479) );
  OR2X1_RVT U4012 ( .A1(n12545), .A2(n3275), .Y(n3314) );
  OR2X1_RVT U4013 ( .A1(n12736), .A2(n3548), .Y(n4055) );
  OR2X1_RVT U4014 ( .A1(n12569), .A2(n3582), .Y(n3548) );
  OR2X1_RVT U4015 ( .A1(n12728), .A2(n12723), .Y(n3582) );
  OR2X1_RVT U4016 ( .A1(n12726), .A2(n12561), .Y(n3258) );
  AND2X1_RVT U4017 ( .A1(n4057), .A2(n4058), .Y(n3452) );
  OR2X1_RVT U4018 ( .A1(n3334), .A2(n3320), .Y(n4058) );
  OR2X1_RVT U4019 ( .A1(n12735), .A2(n3292), .Y(n3320) );
  AND2X1_RVT U4020 ( .A1(n3319), .A2(n3283), .Y(n3372) );
  OR2X1_RVT U4021 ( .A1(n12556), .A2(n3386), .Y(n3334) );
  OR2X1_RVT U4022 ( .A1(n12724), .A2(n3423), .Y(n3386) );
  OR2X1_RVT U4023 ( .A1(n4059), .A2(n3377), .Y(n4057) );
  OR2X1_RVT U4024 ( .A1(n12550), .A2(n254), .Y(n3377) );
  AND2X1_RVT U4025 ( .A1(n12737), .A2(n12543), .Y(n3640) );
  OR2X1_RVT U4026 ( .A1(n12549), .A2(n3480), .Y(n4059) );
  OR2X1_RVT U4027 ( .A1(n12733), .A2(n12566), .Y(n3480) );
  AND2X1_RVT U4028 ( .A1(n4060), .A2(n4061), .Y(n4052) );
  OR2X1_RVT U4029 ( .A1(n3300), .A2(n3633), .Y(n4061) );
  OR2X1_RVT U4030 ( .A1(n12551), .A2(n3340), .Y(n3633) );
  OR2X1_RVT U4031 ( .A1(n12566), .A2(n3417), .Y(n3340) );
  OR2X1_RVT U4032 ( .A1(n12546), .A2(n12549), .Y(n3417) );
  OR2X1_RVT U4033 ( .A1(n12730), .A2(n12728), .Y(n3279) );
  OR2X1_RVT U4034 ( .A1(n12738), .A2(n12732), .Y(n3300) );
  XOR2X1_RVT U4035 ( .A1(key[28]), .A2(state[28]), .Y(n3275) );
  OR2X1_RVT U4036 ( .A1(n3292), .A2(n3421), .Y(n4060) );
  OR2X1_RVT U4037 ( .A1(n3523), .A2(n3714), .Y(n3421) );
  OR2X1_RVT U4038 ( .A1(n12553), .A2(n3321), .Y(n3714) );
  OR2X1_RVT U4039 ( .A1(n12731), .A2(n3423), .Y(n3321) );
  XOR2X1_RVT U4040 ( .A1(key[26]), .A2(state[26]), .Y(n3423) );
  XOR2X1_RVT U4041 ( .A1(key[27]), .A2(state[27]), .Y(n3357) );
  OR2X1_RVT U4042 ( .A1(n12736), .A2(n12551), .Y(n3297) );
  XOR2X1_RVT U4043 ( .A1(key[29]), .A2(state[29]), .Y(n3283) );
  XOR2X1_RVT U4044 ( .A1(key[30]), .A2(state[30]), .Y(n3319) );
  OR2X1_RVT U4045 ( .A1(n12726), .A2(n12549), .Y(n3523) );
  XOR2X1_RVT U4046 ( .A1(key[24]), .A2(state[24]), .Y(n3298) );
  XOR2X1_RVT U4047 ( .A1(key[25]), .A2(state[25]), .Y(n3408) );
  XOR2X1_RVT U4048 ( .A1(key[31]), .A2(state[31]), .Y(n3292) );
  AND4X1_RVT U4049 ( .A1(n4063), .A2(n4064), .A3(n4065), .A4(n4066), .Y(n4062)
         );
  AND4X1_RVT U4050 ( .A1(n4067), .A2(n4068), .A3(n4069), .A4(n4070), .Y(n4066)
         );
  AND4X1_RVT U4051 ( .A1(n4071), .A2(n4072), .A3(n4073), .A4(n4074), .Y(n4070)
         );
  OR2X1_RVT U4052 ( .A1(n12537), .A2(n4076), .Y(n4069) );
  OR2X1_RVT U4053 ( .A1(n4077), .A2(n4078), .Y(n4067) );
  OR2X1_RVT U4054 ( .A1(n12720), .A2(n4079), .Y(n4078) );
  AND4X1_RVT U4055 ( .A1(n4080), .A2(n4081), .A3(n4082), .A4(n4083), .Y(n4065)
         );
  OR2X1_RVT U4056 ( .A1(n4084), .A2(n12718), .Y(n4083) );
  AND2X1_RVT U4057 ( .A1(n4085), .A2(n4086), .Y(n4084) );
  AND2X1_RVT U4058 ( .A1(n4087), .A2(n4088), .Y(n4082) );
  OR2X1_RVT U4059 ( .A1(n4089), .A2(n276), .Y(n4088) );
  AND2X1_RVT U4060 ( .A1(n4090), .A2(n4091), .Y(n4089) );
  OR2X1_RVT U4061 ( .A1(n12528), .A2(n4093), .Y(n4091) );
  OR2X1_RVT U4062 ( .A1(n4079), .A2(n4094), .Y(n4090) );
  OR2X1_RVT U4063 ( .A1(n4095), .A2(n12534), .Y(n4087) );
  AND2X1_RVT U4064 ( .A1(n4097), .A2(n4098), .Y(n4095) );
  OR2X1_RVT U4065 ( .A1(n4099), .A2(n4100), .Y(n4081) );
  AND2X1_RVT U4066 ( .A1(n4101), .A2(n4102), .Y(n4099) );
  OR2X1_RVT U4067 ( .A1(n12529), .A2(n4103), .Y(n4102) );
  AND2X1_RVT U4068 ( .A1(n4104), .A2(n4105), .Y(n4101) );
  AND2X1_RVT U4069 ( .A1(n4106), .A2(n4107), .Y(n4080) );
  OR2X1_RVT U4070 ( .A1(n4108), .A2(n12511), .Y(n4107) );
  AND2X1_RVT U4071 ( .A1(n4110), .A2(n4111), .Y(n4108) );
  OR2X1_RVT U4072 ( .A1(n4112), .A2(n4113), .Y(n4111) );
  OR2X1_RVT U4073 ( .A1(n12520), .A2(n12515), .Y(n4113) );
  OR2X1_RVT U4074 ( .A1(n4116), .A2(n4117), .Y(n4106) );
  AND2X1_RVT U4075 ( .A1(n4118), .A2(n4119), .Y(n4116) );
  AND2X1_RVT U4076 ( .A1(n4120), .A2(n4121), .Y(n4118) );
  AND4X1_RVT U4077 ( .A1(n4122), .A2(n4123), .A3(n4124), .A4(n4125), .Y(n4064)
         );
  AND4X1_RVT U4078 ( .A1(n4126), .A2(n4127), .A3(n4128), .A4(n4129), .Y(n4125)
         );
  OR2X1_RVT U4079 ( .A1(n4130), .A2(n12540), .Y(n4129) );
  AND4X1_RVT U4080 ( .A1(n4132), .A2(n4133), .A3(n4134), .A4(n4135), .Y(n4130)
         );
  OR2X1_RVT U4081 ( .A1(n4136), .A2(n4103), .Y(n4135) );
  OR2X1_RVT U4082 ( .A1(n4137), .A2(n12526), .Y(n4134) );
  OR2X1_RVT U4083 ( .A1(n4139), .A2(n12517), .Y(n4128) );
  AND4X1_RVT U4084 ( .A1(n4140), .A2(n4141), .A3(n4142), .A4(n4143), .Y(n4139)
         );
  OR2X1_RVT U4085 ( .A1(n4144), .A2(n4145), .Y(n4143) );
  OR2X1_RVT U4086 ( .A1(n12534), .A2(n12529), .Y(n4145) );
  AND2X1_RVT U4087 ( .A1(n4146), .A2(n4147), .Y(n4142) );
  OR2X1_RVT U4088 ( .A1(n12722), .A2(n4148), .Y(n4141) );
  OR2X1_RVT U4089 ( .A1(n4149), .A2(n4150), .Y(n4140) );
  AND2X1_RVT U4090 ( .A1(n4151), .A2(n4152), .Y(n4149) );
  OR2X1_RVT U4091 ( .A1(n12534), .A2(n4153), .Y(n4152) );
  OR2X1_RVT U4092 ( .A1(n4086), .A2(n4154), .Y(n4127) );
  OR2X1_RVT U4093 ( .A1(n4153), .A2(n4155), .Y(n4126) );
  OR2X1_RVT U4094 ( .A1(n4156), .A2(n4157), .Y(n4124) );
  OR2X1_RVT U4095 ( .A1(n4158), .A2(n4151), .Y(n4123) );
  OR2X1_RVT U4096 ( .A1(n4159), .A2(n4160), .Y(n4122) );
  AND4X1_RVT U4097 ( .A1(n4161), .A2(n4162), .A3(n4163), .A4(n4164), .Y(n4063)
         );
  AND2X1_RVT U4098 ( .A1(n4165), .A2(n4166), .Y(n4164) );
  OR2X1_RVT U4099 ( .A1(n4150), .A2(n4167), .Y(n4166) );
  AND2X1_RVT U4100 ( .A1(n4168), .A2(n4169), .Y(n4165) );
  OR2X1_RVT U4101 ( .A1(n4170), .A2(n4093), .Y(n4169) );
  OR2X1_RVT U4102 ( .A1(n4094), .A2(n4171), .Y(n4168) );
  OR2X1_RVT U4103 ( .A1(n274), .A2(n4172), .Y(n4163) );
  OR2X1_RVT U4104 ( .A1(n4173), .A2(n12524), .Y(n4162) );
  OR2X1_RVT U4105 ( .A1(n12527), .A2(n4175), .Y(n4161) );
  AND4X1_RVT U4106 ( .A1(n4177), .A2(n4178), .A3(n4179), .A4(n4180), .Y(n4176)
         );
  AND4X1_RVT U4107 ( .A1(n4181), .A2(n4072), .A3(n4182), .A4(n4183), .Y(n4180)
         );
  AND4X1_RVT U4108 ( .A1(n4184), .A2(n4185), .A3(n4186), .A4(n4187), .Y(n4183)
         );
  OR2X1_RVT U4109 ( .A1(n4093), .A2(n4188), .Y(n4187) );
  OR2X1_RVT U4110 ( .A1(n4189), .A2(n12539), .Y(n4188) );
  OR2X1_RVT U4111 ( .A1(n4094), .A2(n4190), .Y(n4186) );
  OR2X1_RVT U4112 ( .A1(n274), .A2(n12523), .Y(n4190) );
  OR2X1_RVT U4113 ( .A1(n4191), .A2(n4137), .Y(n4185) );
  AND2X1_RVT U4114 ( .A1(n4148), .A2(n4192), .Y(n4191) );
  OR2X1_RVT U4115 ( .A1(n4193), .A2(n4194), .Y(n4184) );
  AND2X1_RVT U4116 ( .A1(n4195), .A2(n4196), .Y(n4193) );
  AND2X1_RVT U4117 ( .A1(n4197), .A2(n4198), .Y(n4182) );
  OR2X1_RVT U4118 ( .A1(n4144), .A2(n4199), .Y(n4198) );
  OR2X1_RVT U4119 ( .A1(n4200), .A2(n12720), .Y(n4199) );
  OR2X1_RVT U4120 ( .A1(n4201), .A2(n4202), .Y(n4197) );
  OR2X1_RVT U4121 ( .A1(n4203), .A2(n12528), .Y(n4202) );
  OR2X1_RVT U4122 ( .A1(n4079), .A2(n4204), .Y(n4072) );
  AND4X1_RVT U4123 ( .A1(n4205), .A2(n4206), .A3(n4207), .A4(n4208), .Y(n4179)
         );
  AND4X1_RVT U4124 ( .A1(n4209), .A2(n4210), .A3(n4211), .A4(n4212), .Y(n4208)
         );
  OR2X1_RVT U4125 ( .A1(n4213), .A2(n12542), .Y(n4212) );
  AND2X1_RVT U4126 ( .A1(n4215), .A2(n4216), .Y(n4213) );
  OR2X1_RVT U4127 ( .A1(n12511), .A2(n4094), .Y(n4216) );
  OR2X1_RVT U4128 ( .A1(n4217), .A2(n4096), .Y(n4211) );
  AND2X1_RVT U4129 ( .A1(n4218), .A2(n4219), .Y(n4217) );
  OR2X1_RVT U4130 ( .A1(n4220), .A2(n12719), .Y(n4210) );
  AND2X1_RVT U4131 ( .A1(n4221), .A2(n4222), .Y(n4220) );
  OR2X1_RVT U4132 ( .A1(n4223), .A2(n4172), .Y(n4222) );
  AND2X1_RVT U4133 ( .A1(n12542), .A2(n12526), .Y(n4223) );
  OR2X1_RVT U4134 ( .A1(n4224), .A2(n12512), .Y(n4209) );
  AND2X1_RVT U4135 ( .A1(n4226), .A2(n4227), .Y(n4224) );
  OR2X1_RVT U4136 ( .A1(n4228), .A2(n12518), .Y(n4207) );
  AND2X1_RVT U4137 ( .A1(n4229), .A2(n4230), .Y(n4228) );
  OR2X1_RVT U4138 ( .A1(n12526), .A2(n4231), .Y(n4230) );
  AND2X1_RVT U4139 ( .A1(n4232), .A2(n4233), .Y(n4229) );
  OR2X1_RVT U4140 ( .A1(n4234), .A2(n4235), .Y(n4232) );
  OR2X1_RVT U4141 ( .A1(n4079), .A2(n4150), .Y(n4235) );
  OR2X1_RVT U4142 ( .A1(n4236), .A2(n12716), .Y(n4206) );
  AND2X1_RVT U4143 ( .A1(n4237), .A2(n4238), .Y(n4236) );
  OR2X1_RVT U4144 ( .A1(n4239), .A2(n4240), .Y(n4205) );
  AND2X1_RVT U4145 ( .A1(n4241), .A2(n4242), .Y(n4239) );
  AND2X1_RVT U4146 ( .A1(n4243), .A2(n4244), .Y(n4241) );
  OR2X1_RVT U4147 ( .A1(n276), .A2(n4172), .Y(n4244) );
  OR2X1_RVT U4148 ( .A1(n12536), .A2(n4137), .Y(n4243) );
  AND4X1_RVT U4149 ( .A1(n4245), .A2(n4246), .A3(n4247), .A4(n4248), .Y(n4178)
         );
  AND4X1_RVT U4150 ( .A1(n4249), .A2(n4250), .A3(n4251), .A4(n4252), .Y(n4248)
         );
  OR2X1_RVT U4151 ( .A1(n4172), .A2(n4171), .Y(n4252) );
  OR2X1_RVT U4152 ( .A1(n4103), .A2(n4253), .Y(n4251) );
  OR2X1_RVT U4153 ( .A1(n4136), .A2(n4254), .Y(n4250) );
  OR2X1_RVT U4154 ( .A1(n4079), .A2(n4255), .Y(n4249) );
  AND2X1_RVT U4155 ( .A1(n4256), .A2(n4257), .Y(n4247) );
  OR2X1_RVT U4156 ( .A1(n12537), .A2(n4258), .Y(n4257) );
  OR2X1_RVT U4157 ( .A1(n12516), .A2(n4155), .Y(n4256) );
  OR2X1_RVT U4158 ( .A1(n4259), .A2(n4114), .Y(n4246) );
  AND4X1_RVT U4159 ( .A1(n4260), .A2(n4261), .A3(n4262), .A4(n4263), .Y(n4259)
         );
  OR2X1_RVT U4160 ( .A1(n4264), .A2(n4079), .Y(n4262) );
  OR2X1_RVT U4161 ( .A1(n12708), .A2(n4265), .Y(n4261) );
  OR2X1_RVT U4162 ( .A1(n4266), .A2(n12716), .Y(n4260) );
  AND2X1_RVT U4163 ( .A1(n4157), .A2(n4267), .Y(n4266) );
  OR2X1_RVT U4164 ( .A1(n4159), .A2(n4268), .Y(n4245) );
  AND4X1_RVT U4165 ( .A1(n4269), .A2(n4270), .A3(n4271), .A4(n4272), .Y(n4177)
         );
  AND4X1_RVT U4166 ( .A1(n4273), .A2(n4274), .A3(n4275), .A4(n4276), .Y(n4272)
         );
  OR2X1_RVT U4167 ( .A1(n12712), .A2(n4277), .Y(n4276) );
  OR2X1_RVT U4168 ( .A1(n12713), .A2(n4278), .Y(n4275) );
  OR2X1_RVT U4169 ( .A1(n12710), .A2(n4279), .Y(n4274) );
  OR2X1_RVT U4170 ( .A1(n12510), .A2(n4280), .Y(n4273) );
  OR2X1_RVT U4171 ( .A1(n4281), .A2(n12517), .Y(n4270) );
  AND4X1_RVT U4172 ( .A1(n4283), .A2(n4284), .A3(n4285), .A4(n4286), .Y(n4282)
         );
  AND4X1_RVT U4173 ( .A1(n4287), .A2(n4288), .A3(n4289), .A4(n4290), .Y(n4286)
         );
  AND4X1_RVT U4174 ( .A1(n4291), .A2(n4068), .A3(n4238), .A4(n4292), .Y(n4290)
         );
  OR2X1_RVT U4175 ( .A1(n4293), .A2(n12707), .Y(n4068) );
  AND2X1_RVT U4176 ( .A1(n4294), .A2(n4295), .Y(n4293) );
  OR2X1_RVT U4177 ( .A1(n4112), .A2(n4296), .Y(n4295) );
  OR2X1_RVT U4178 ( .A1(n4297), .A2(n4194), .Y(n4294) );
  OR2X1_RVT U4179 ( .A1(n4298), .A2(n4153), .Y(n4291) );
  AND2X1_RVT U4180 ( .A1(n4299), .A2(n4300), .Y(n4298) );
  OR2X1_RVT U4181 ( .A1(n12712), .A2(n4137), .Y(n4300) );
  OR2X1_RVT U4182 ( .A1(n4301), .A2(n4096), .Y(n4289) );
  AND2X1_RVT U4183 ( .A1(n4302), .A2(n4303), .Y(n4301) );
  OR2X1_RVT U4184 ( .A1(n4304), .A2(n12718), .Y(n4303) );
  AND2X1_RVT U4185 ( .A1(n4144), .A2(n4305), .Y(n4304) );
  OR2X1_RVT U4186 ( .A1(n4306), .A2(n12537), .Y(n4288) );
  AND2X1_RVT U4187 ( .A1(n4307), .A2(n4308), .Y(n4306) );
  OR2X1_RVT U4188 ( .A1(n4137), .A2(n4103), .Y(n4308) );
  OR2X1_RVT U4189 ( .A1(n4309), .A2(n12520), .Y(n4287) );
  AND2X1_RVT U4190 ( .A1(n4221), .A2(n4310), .Y(n4309) );
  OR2X1_RVT U4191 ( .A1(n4150), .A2(n4311), .Y(n4221) );
  AND4X1_RVT U4192 ( .A1(n4312), .A2(n4313), .A3(n4314), .A4(n4315), .Y(n4285)
         );
  OR2X1_RVT U4193 ( .A1(n4316), .A2(n12527), .Y(n4315) );
  AND2X1_RVT U4194 ( .A1(n4317), .A2(n4318), .Y(n4316) );
  OR2X1_RVT U4195 ( .A1(n4194), .A2(n4094), .Y(n4318) );
  AND2X1_RVT U4196 ( .A1(n4319), .A2(n4320), .Y(n4317) );
  OR2X1_RVT U4197 ( .A1(n4234), .A2(n4296), .Y(n4319) );
  AND2X1_RVT U4198 ( .A1(n4321), .A2(n4322), .Y(n4314) );
  OR2X1_RVT U4199 ( .A1(n4323), .A2(n4225), .Y(n4322) );
  AND2X1_RVT U4200 ( .A1(n4324), .A2(n4133), .Y(n4323) );
  OR2X1_RVT U4201 ( .A1(n4079), .A2(n4194), .Y(n4133) );
  OR2X1_RVT U4202 ( .A1(n4325), .A2(n276), .Y(n4321) );
  AND2X1_RVT U4203 ( .A1(n4326), .A2(n4327), .Y(n4325) );
  OR2X1_RVT U4204 ( .A1(n4328), .A2(n12529), .Y(n4327) );
  AND2X1_RVT U4205 ( .A1(n4329), .A2(n4330), .Y(n4328) );
  OR2X1_RVT U4206 ( .A1(n12524), .A2(n4144), .Y(n4330) );
  OR2X1_RVT U4207 ( .A1(n12722), .A2(n12526), .Y(n4329) );
  AND2X1_RVT U4208 ( .A1(n4195), .A2(n4305), .Y(n4326) );
  OR2X1_RVT U4209 ( .A1(n4225), .A2(n4331), .Y(n4195) );
  OR2X1_RVT U4210 ( .A1(n12717), .A2(n12713), .Y(n4331) );
  OR2X1_RVT U4211 ( .A1(n4332), .A2(n4214), .Y(n4313) );
  AND4X1_RVT U4212 ( .A1(n4173), .A2(n4333), .A3(n4334), .A4(n4335), .Y(n4332)
         );
  OR2X1_RVT U4213 ( .A1(n12528), .A2(n4194), .Y(n4335) );
  AND2X1_RVT U4214 ( .A1(n4336), .A2(n4337), .Y(n4334) );
  OR2X1_RVT U4215 ( .A1(n12722), .A2(n12537), .Y(n4333) );
  AND2X1_RVT U4216 ( .A1(n4338), .A2(n4339), .Y(n4173) );
  OR2X1_RVT U4217 ( .A1(n4340), .A2(n274), .Y(n4339) );
  OR2X1_RVT U4218 ( .A1(n4137), .A2(n12707), .Y(n4338) );
  AND2X1_RVT U4219 ( .A1(n4341), .A2(n4342), .Y(n4312) );
  OR2X1_RVT U4220 ( .A1(n4343), .A2(n12709), .Y(n4342) );
  AND2X1_RVT U4221 ( .A1(n4344), .A2(n4345), .Y(n4343) );
  OR2X1_RVT U4222 ( .A1(n4346), .A2(n12531), .Y(n4345) );
  AND2X1_RVT U4223 ( .A1(n4347), .A2(n4348), .Y(n4346) );
  AND2X1_RVT U4224 ( .A1(n4349), .A2(n4350), .Y(n4344) );
  OR2X1_RVT U4225 ( .A1(n4351), .A2(n12540), .Y(n4341) );
  AND4X1_RVT U4226 ( .A1(n4352), .A2(n4353), .A3(n4354), .A4(n4355), .Y(n4351)
         );
  OR2X1_RVT U4227 ( .A1(n12721), .A2(n4356), .Y(n4354) );
  OR2X1_RVT U4228 ( .A1(n274), .A2(n4151), .Y(n4353) );
  OR2X1_RVT U4229 ( .A1(n4240), .A2(n4194), .Y(n4352) );
  AND4X1_RVT U4230 ( .A1(n4357), .A2(n4358), .A3(n4359), .A4(n4360), .Y(n4284)
         );
  AND2X1_RVT U4231 ( .A1(n4361), .A2(n4204), .Y(n4360) );
  OR2X1_RVT U4232 ( .A1(n12515), .A2(n4170), .Y(n4204) );
  AND2X1_RVT U4233 ( .A1(n4362), .A2(n4363), .Y(n4361) );
  OR2X1_RVT U4234 ( .A1(n4364), .A2(n4119), .Y(n4363) );
  OR2X1_RVT U4235 ( .A1(n4171), .A2(n4231), .Y(n4362) );
  OR2X1_RVT U4236 ( .A1(n274), .A2(n4365), .Y(n4359) );
  OR2X1_RVT U4237 ( .A1(n12720), .A2(n4366), .Y(n4358) );
  OR2X1_RVT U4238 ( .A1(n4240), .A2(n4367), .Y(n4357) );
  AND4X1_RVT U4239 ( .A1(n4368), .A2(n4369), .A3(n4370), .A4(n4371), .Y(n4283)
         );
  AND2X1_RVT U4240 ( .A1(n4372), .A2(n4373), .Y(n4371) );
  OR2X1_RVT U4241 ( .A1(n12510), .A2(n4374), .Y(n4373) );
  AND2X1_RVT U4242 ( .A1(n4375), .A2(n4376), .Y(n4372) );
  OR2X1_RVT U4243 ( .A1(n4136), .A2(n4146), .Y(n4376) );
  OR2X1_RVT U4244 ( .A1(n12531), .A2(n4196), .Y(n4146) );
  OR2X1_RVT U4245 ( .A1(n12517), .A2(n4377), .Y(n4375) );
  OR2X1_RVT U4246 ( .A1(n4117), .A2(n4110), .Y(n4370) );
  OR2X1_RVT U4247 ( .A1(n4203), .A2(n4378), .Y(n4110) );
  OR2X1_RVT U4248 ( .A1(n12716), .A2(n4379), .Y(n4369) );
  OR2X1_RVT U4249 ( .A1(n12529), .A2(n4237), .Y(n4368) );
  OR2X1_RVT U4250 ( .A1(n12707), .A2(n4299), .Y(n4237) );
  AND4X1_RVT U4251 ( .A1(n4381), .A2(n4382), .A3(n4383), .A4(n4384), .Y(n4380)
         );
  AND4X1_RVT U4252 ( .A1(n4385), .A2(n4386), .A3(n4387), .A4(n4388), .Y(n4384)
         );
  OR2X1_RVT U4253 ( .A1(n284), .A2(n4389), .Y(n4388) );
  OR2X1_RVT U4254 ( .A1(n4390), .A2(n12542), .Y(n4389) );
  AND2X1_RVT U4255 ( .A1(n12531), .A2(n4156), .Y(n4390) );
  AND2X1_RVT U4256 ( .A1(n4071), .A2(n4391), .Y(n4387) );
  OR2X1_RVT U4257 ( .A1(n12520), .A2(n4392), .Y(n4071) );
  OR2X1_RVT U4258 ( .A1(n284), .A2(n4150), .Y(n4392) );
  OR2X1_RVT U4259 ( .A1(n4393), .A2(n4079), .Y(n4386) );
  AND2X1_RVT U4260 ( .A1(n4394), .A2(n4395), .Y(n4393) );
  AND2X1_RVT U4261 ( .A1(n4396), .A2(n4397), .Y(n4385) );
  OR2X1_RVT U4262 ( .A1(n4398), .A2(n4399), .Y(n4397) );
  AND2X1_RVT U4263 ( .A1(n4400), .A2(n4160), .Y(n4398) );
  OR2X1_RVT U4264 ( .A1(n4401), .A2(n4151), .Y(n4396) );
  AND2X1_RVT U4265 ( .A1(n4336), .A2(n4170), .Y(n4401) );
  OR2X1_RVT U4266 ( .A1(n12518), .A2(n4402), .Y(n4336) );
  OR2X1_RVT U4267 ( .A1(n12722), .A2(n12528), .Y(n4402) );
  AND4X1_RVT U4268 ( .A1(n4403), .A2(n4404), .A3(n4405), .A4(n4406), .Y(n4383)
         );
  OR2X1_RVT U4269 ( .A1(n4407), .A2(n12712), .Y(n4406) );
  AND2X1_RVT U4270 ( .A1(n4219), .A2(n4408), .Y(n4407) );
  OR2X1_RVT U4271 ( .A1(n12720), .A2(n4264), .Y(n4219) );
  AND2X1_RVT U4272 ( .A1(n4409), .A2(n4410), .Y(n4405) );
  OR2X1_RVT U4273 ( .A1(n4411), .A2(n12710), .Y(n4410) );
  AND2X1_RVT U4274 ( .A1(n4412), .A2(n4413), .Y(n4411) );
  OR2X1_RVT U4275 ( .A1(n4114), .A2(n4356), .Y(n4413) );
  OR2X1_RVT U4276 ( .A1(n4414), .A2(n12708), .Y(n4409) );
  AND2X1_RVT U4277 ( .A1(n4415), .A2(n4416), .Y(n4414) );
  OR2X1_RVT U4278 ( .A1(n4417), .A2(n12531), .Y(n4404) );
  AND2X1_RVT U4279 ( .A1(n4418), .A2(n4419), .Y(n4417) );
  AND2X1_RVT U4280 ( .A1(n4420), .A2(n4421), .Y(n4418) );
  AND2X1_RVT U4281 ( .A1(n4422), .A2(n4423), .Y(n4403) );
  OR2X1_RVT U4282 ( .A1(n4424), .A2(n4340), .Y(n4423) );
  AND2X1_RVT U4283 ( .A1(n4425), .A2(n4171), .Y(n4424) );
  AND2X1_RVT U4284 ( .A1(n4426), .A2(n4427), .Y(n4425) );
  OR2X1_RVT U4285 ( .A1(n4428), .A2(n12534), .Y(n4422) );
  AND2X1_RVT U4286 ( .A1(n4429), .A2(n4430), .Y(n4428) );
  OR2X1_RVT U4287 ( .A1(n12719), .A2(n12536), .Y(n4430) );
  AND2X1_RVT U4288 ( .A1(n4160), .A2(n4431), .Y(n4429) );
  AND4X1_RVT U4289 ( .A1(n4432), .A2(n4433), .A3(n4434), .A4(n4435), .Y(n4382)
         );
  AND2X1_RVT U4290 ( .A1(n4436), .A2(n4437), .Y(n4435) );
  OR2X1_RVT U4291 ( .A1(n4153), .A2(n4227), .Y(n4437) );
  OR2X1_RVT U4292 ( .A1(n12714), .A2(n4160), .Y(n4227) );
  AND2X1_RVT U4293 ( .A1(n4438), .A2(n4439), .Y(n4436) );
  OR2X1_RVT U4294 ( .A1(n4305), .A2(n4119), .Y(n4439) );
  OR2X1_RVT U4295 ( .A1(n12721), .A2(n12527), .Y(n4119) );
  OR2X1_RVT U4296 ( .A1(n4203), .A2(n4253), .Y(n4438) );
  OR2X1_RVT U4297 ( .A1(n12709), .A2(n4440), .Y(n4253) );
  OR2X1_RVT U4298 ( .A1(n4441), .A2(n12510), .Y(n4434) );
  AND4X1_RVT U4299 ( .A1(n4442), .A2(n4443), .A3(n4444), .A4(n4445), .Y(n4441)
         );
  OR2X1_RVT U4300 ( .A1(n4378), .A2(n4151), .Y(n4444) );
  OR2X1_RVT U4301 ( .A1(n4446), .A2(n4148), .Y(n4443) );
  OR2X1_RVT U4302 ( .A1(n12718), .A2(n4103), .Y(n4442) );
  OR2X1_RVT U4303 ( .A1(n4447), .A2(n12511), .Y(n4433) );
  AND2X1_RVT U4304 ( .A1(n4448), .A2(n4449), .Y(n4447) );
  OR2X1_RVT U4305 ( .A1(n4378), .A2(n4103), .Y(n4449) );
  AND2X1_RVT U4306 ( .A1(n4450), .A2(n4379), .Y(n4448) );
  OR2X1_RVT U4307 ( .A1(n4151), .A2(n4451), .Y(n4379) );
  OR2X1_RVT U4308 ( .A1(n12709), .A2(n12721), .Y(n4451) );
  OR2X1_RVT U4309 ( .A1(n4452), .A2(n12518), .Y(n4432) );
  AND4X1_RVT U4310 ( .A1(n4453), .A2(n4366), .A3(n4175), .A4(n4147), .Y(n4452)
         );
  OR2X1_RVT U4311 ( .A1(n4172), .A2(n4454), .Y(n4147) );
  OR2X1_RVT U4312 ( .A1(n12711), .A2(n4109), .Y(n4454) );
  OR2X1_RVT U4313 ( .A1(n4234), .A2(n4268), .Y(n4175) );
  OR2X1_RVT U4314 ( .A1(n4153), .A2(n4455), .Y(n4366) );
  OR2X1_RVT U4315 ( .A1(n12542), .A2(n12511), .Y(n4455) );
  OR2X1_RVT U4316 ( .A1(n4112), .A2(n4456), .Y(n4453) );
  OR2X1_RVT U4317 ( .A1(n4457), .A2(n12516), .Y(n4456) );
  AND4X1_RVT U4318 ( .A1(n4458), .A2(n4459), .A3(n4460), .A4(n4461), .Y(n4381)
         );
  AND2X1_RVT U4319 ( .A1(n4462), .A2(n4463), .Y(n4461) );
  AND2X1_RVT U4320 ( .A1(n4464), .A2(n4465), .Y(n4462) );
  OR2X1_RVT U4321 ( .A1(n4144), .A2(n4419), .Y(n4465) );
  OR2X1_RVT U4322 ( .A1(n4156), .A2(n4466), .Y(n4419) );
  OR2X1_RVT U4323 ( .A1(n12710), .A2(n12712), .Y(n4466) );
  OR2X1_RVT U4324 ( .A1(n12717), .A2(n4467), .Y(n4464) );
  OR2X1_RVT U4325 ( .A1(n12527), .A2(n4468), .Y(n4460) );
  OR2X1_RVT U4326 ( .A1(n12720), .A2(n4469), .Y(n4459) );
  OR2X1_RVT U4327 ( .A1(n4156), .A2(n4470), .Y(n4458) );
  AND4X1_RVT U4328 ( .A1(n4472), .A2(n4473), .A3(n4474), .A4(n4475), .Y(n4471)
         );
  AND4X1_RVT U4329 ( .A1(n4476), .A2(n4477), .A3(n4478), .A4(n4479), .Y(n4475)
         );
  AND4X1_RVT U4330 ( .A1(n4480), .A2(n4481), .A3(n4073), .A4(n4482), .Y(n4479)
         );
  OR2X1_RVT U4331 ( .A1(n4214), .A2(n4483), .Y(n4073) );
  OR2X1_RVT U4332 ( .A1(n4305), .A2(n276), .Y(n4483) );
  OR2X1_RVT U4333 ( .A1(n4077), .A2(n4484), .Y(n4481) );
  OR2X1_RVT U4334 ( .A1(n12715), .A2(n12718), .Y(n4484) );
  OR2X1_RVT U4335 ( .A1(n4340), .A2(n4485), .Y(n4480) );
  OR2X1_RVT U4336 ( .A1(n4486), .A2(n4114), .Y(n4485) );
  AND2X1_RVT U4337 ( .A1(n12531), .A2(n4214), .Y(n4486) );
  OR2X1_RVT U4338 ( .A1(n4487), .A2(n12537), .Y(n4478) );
  AND2X1_RVT U4339 ( .A1(n4355), .A2(n4427), .Y(n4487) );
  OR2X1_RVT U4340 ( .A1(n276), .A2(n4488), .Y(n4427) );
  OR2X1_RVT U4341 ( .A1(n12510), .A2(n12714), .Y(n4488) );
  OR2X1_RVT U4342 ( .A1(n4144), .A2(n4489), .Y(n4355) );
  OR2X1_RVT U4343 ( .A1(n12712), .A2(n4136), .Y(n4489) );
  OR2X1_RVT U4344 ( .A1(n4490), .A2(n4094), .Y(n4477) );
  AND2X1_RVT U4345 ( .A1(n4491), .A2(n4299), .Y(n4490) );
  OR2X1_RVT U4346 ( .A1(n4200), .A2(n4194), .Y(n4476) );
  AND4X1_RVT U4347 ( .A1(n4492), .A2(n4493), .A3(n4494), .A4(n4495), .Y(n4474)
         );
  AND2X1_RVT U4348 ( .A1(n4496), .A2(n4497), .Y(n4495) );
  OR2X1_RVT U4349 ( .A1(n4498), .A2(n12531), .Y(n4497) );
  AND2X1_RVT U4350 ( .A1(n4499), .A2(n4167), .Y(n4498) );
  AND2X1_RVT U4351 ( .A1(n4500), .A2(n4501), .Y(n4496) );
  OR2X1_RVT U4352 ( .A1(n4502), .A2(n4150), .Y(n4501) );
  AND2X1_RVT U4353 ( .A1(n4121), .A2(n4093), .Y(n4502) );
  OR2X1_RVT U4354 ( .A1(n12720), .A2(n4192), .Y(n4121) );
  OR2X1_RVT U4355 ( .A1(n4503), .A2(n4203), .Y(n4500) );
  AND2X1_RVT U4356 ( .A1(n4395), .A2(n4504), .Y(n4503) );
  OR2X1_RVT U4357 ( .A1(n12721), .A2(n4231), .Y(n4395) );
  OR2X1_RVT U4358 ( .A1(n4505), .A2(n12712), .Y(n4494) );
  AND2X1_RVT U4359 ( .A1(n4098), .A2(n4506), .Y(n4505) );
  OR2X1_RVT U4360 ( .A1(n4234), .A2(n4158), .Y(n4506) );
  OR2X1_RVT U4361 ( .A1(n4137), .A2(n4340), .Y(n4098) );
  OR2X1_RVT U4362 ( .A1(n4507), .A2(n274), .Y(n4493) );
  AND2X1_RVT U4363 ( .A1(n4148), .A2(n4508), .Y(n4507) );
  OR2X1_RVT U4364 ( .A1(n4509), .A2(n12515), .Y(n4508) );
  AND2X1_RVT U4365 ( .A1(n4510), .A2(n4511), .Y(n4509) );
  OR2X1_RVT U4366 ( .A1(n12713), .A2(n4131), .Y(n4511) );
  OR2X1_RVT U4367 ( .A1(n12542), .A2(n4234), .Y(n4148) );
  OR2X1_RVT U4368 ( .A1(n4512), .A2(n4218), .Y(n4492) );
  AND2X1_RVT U4369 ( .A1(n4151), .A2(n4196), .Y(n4512) );
  OR2X1_RVT U4370 ( .A1(n12709), .A2(n4079), .Y(n4196) );
  AND4X1_RVT U4371 ( .A1(n4513), .A2(n4514), .A3(n4515), .A4(n4516), .Y(n4473)
         );
  AND4X1_RVT U4372 ( .A1(n4517), .A2(n4518), .A3(n4519), .A4(n4520), .Y(n4516)
         );
  OR2X1_RVT U4373 ( .A1(n4521), .A2(n12720), .Y(n4520) );
  AND2X1_RVT U4374 ( .A1(n4254), .A2(n4522), .Y(n4521) );
  OR2X1_RVT U4375 ( .A1(n12539), .A2(n4103), .Y(n4522) );
  OR2X1_RVT U4376 ( .A1(n4523), .A2(n4096), .Y(n4519) );
  AND2X1_RVT U4377 ( .A1(n4524), .A2(n4525), .Y(n4523) );
  OR2X1_RVT U4378 ( .A1(n4526), .A2(n4131), .Y(n4525) );
  AND2X1_RVT U4379 ( .A1(n4156), .A2(n4144), .Y(n4526) );
  AND2X1_RVT U4380 ( .A1(n4158), .A2(n4400), .Y(n4524) );
  OR2X1_RVT U4381 ( .A1(n12540), .A2(n4296), .Y(n4400) );
  OR2X1_RVT U4382 ( .A1(n4527), .A2(n12529), .Y(n4518) );
  AND2X1_RVT U4383 ( .A1(n4528), .A2(n4529), .Y(n4527) );
  OR2X1_RVT U4384 ( .A1(n4144), .A2(n4530), .Y(n4529) );
  AND2X1_RVT U4385 ( .A1(n4226), .A2(n4420), .Y(n4528) );
  OR2X1_RVT U4386 ( .A1(n4136), .A2(n4311), .Y(n4420) );
  OR2X1_RVT U4387 ( .A1(n4109), .A2(n4531), .Y(n4226) );
  OR2X1_RVT U4388 ( .A1(n4532), .A2(n4079), .Y(n4517) );
  AND4X1_RVT U4389 ( .A1(n4533), .A2(n4534), .A3(n4535), .A4(n4468), .Y(n4532)
         );
  OR2X1_RVT U4390 ( .A1(n4172), .A2(n4536), .Y(n4468) );
  OR2X1_RVT U4391 ( .A1(n12510), .A2(n4136), .Y(n4536) );
  OR2X1_RVT U4392 ( .A1(n12717), .A2(n4378), .Y(n4534) );
  OR2X1_RVT U4393 ( .A1(n4137), .A2(n4234), .Y(n4533) );
  OR2X1_RVT U4394 ( .A1(n4305), .A2(n4347), .Y(n4515) );
  OR2X1_RVT U4395 ( .A1(n4537), .A2(n12513), .Y(n4514) );
  AND4X1_RVT U4396 ( .A1(n4538), .A2(n4539), .A3(n4181), .A4(n4279), .Y(n4537)
         );
  OR2X1_RVT U4397 ( .A1(n4103), .A2(n4268), .Y(n4279) );
  OR2X1_RVT U4398 ( .A1(n12717), .A2(n274), .Y(n4268) );
  OR2X1_RVT U4399 ( .A1(n4096), .A2(n4160), .Y(n4181) );
  OR2X1_RVT U4400 ( .A1(n12709), .A2(n4531), .Y(n4513) );
  AND4X1_RVT U4401 ( .A1(n4540), .A2(n4541), .A3(n4542), .A4(n4543), .Y(n4472)
         );
  OR2X1_RVT U4402 ( .A1(n12518), .A2(n4544), .Y(n4543) );
  AND2X1_RVT U4403 ( .A1(n4545), .A2(n4546), .Y(n4542) );
  OR2X1_RVT U4404 ( .A1(n12539), .A2(n4299), .Y(n4546) );
  OR2X1_RVT U4405 ( .A1(n4086), .A2(n4160), .Y(n4545) );
  OR2X1_RVT U4406 ( .A1(n276), .A2(n4117), .Y(n4160) );
  OR2X1_RVT U4407 ( .A1(n12542), .A2(n4278), .Y(n4541) );
  OR2X1_RVT U4408 ( .A1(n4153), .A2(n4547), .Y(n4278) );
  AND2X1_RVT U4409 ( .A1(n4548), .A2(n4549), .Y(n4540) );
  OR2X1_RVT U4410 ( .A1(n12511), .A2(n4550), .Y(n4549) );
  OR2X1_RVT U4411 ( .A1(n4156), .A2(n4105), .Y(n4548) );
  OR2X1_RVT U4412 ( .A1(n4079), .A2(n4364), .Y(n4105) );
  AND4X1_RVT U4413 ( .A1(n4552), .A2(n4553), .A3(n4554), .A4(n4555), .Y(n4551)
         );
  AND4X1_RVT U4414 ( .A1(n4556), .A2(n4557), .A3(n4558), .A4(n4559), .Y(n4555)
         );
  AND4X1_RVT U4415 ( .A1(n4292), .A2(n4482), .A3(n4560), .A4(n4561), .Y(n4559)
         );
  OR2X1_RVT U4416 ( .A1(n4562), .A2(n4563), .Y(n4482) );
  OR2X1_RVT U4417 ( .A1(n4077), .A2(n4347), .Y(n4292) );
  OR2X1_RVT U4418 ( .A1(n12718), .A2(n12527), .Y(n4347) );
  AND4X1_RVT U4419 ( .A1(n4550), .A2(n4416), .A3(n4539), .A4(n4074), .Y(n4558)
         );
  OR2X1_RVT U4420 ( .A1(n4564), .A2(n4264), .Y(n4074) );
  OR2X1_RVT U4421 ( .A1(n4079), .A2(n4565), .Y(n4539) );
  OR2X1_RVT U4422 ( .A1(n4112), .A2(n274), .Y(n4416) );
  OR2X1_RVT U4423 ( .A1(n4103), .A2(n4566), .Y(n4550) );
  OR2X1_RVT U4424 ( .A1(n12517), .A2(n12537), .Y(n4566) );
  AND4X1_RVT U4425 ( .A1(n4567), .A2(n4568), .A3(n4569), .A4(n4570), .Y(n4557)
         );
  OR2X1_RVT U4426 ( .A1(n4356), .A2(n4571), .Y(n4570) );
  OR2X1_RVT U4427 ( .A1(n12537), .A2(n4136), .Y(n4571) );
  OR2X1_RVT U4428 ( .A1(n4265), .A2(n4572), .Y(n4569) );
  OR2X1_RVT U4429 ( .A1(n12719), .A2(n4153), .Y(n4572) );
  OR2X1_RVT U4430 ( .A1(n4491), .A2(n4573), .Y(n4568) );
  OR2X1_RVT U4431 ( .A1(n4574), .A2(n4150), .Y(n4573) );
  OR2X1_RVT U4432 ( .A1(n12534), .A2(n4575), .Y(n4567) );
  OR2X1_RVT U4433 ( .A1(n4576), .A2(n12517), .Y(n4575) );
  AND2X1_RVT U4434 ( .A1(n4364), .A2(n4577), .Y(n4576) );
  AND2X1_RVT U4435 ( .A1(n4578), .A2(n4579), .Y(n4556) );
  OR2X1_RVT U4436 ( .A1(n4580), .A2(n4131), .Y(n4579) );
  AND2X1_RVT U4437 ( .A1(n4581), .A2(n4582), .Y(n4580) );
  OR2X1_RVT U4438 ( .A1(n12516), .A2(n4324), .Y(n4582) );
  OR2X1_RVT U4439 ( .A1(n12520), .A2(n4399), .Y(n4581) );
  AND2X1_RVT U4440 ( .A1(n4583), .A2(n4584), .Y(n4578) );
  OR2X1_RVT U4441 ( .A1(n4585), .A2(n4170), .Y(n4584) );
  AND2X1_RVT U4442 ( .A1(n4586), .A2(n4587), .Y(n4585) );
  OR2X1_RVT U4443 ( .A1(n12523), .A2(n284), .Y(n4587) );
  NAND2X1_RVT U4444 ( .A1(n4153), .A2(n12711), .Y(n4586) );
  OR2X1_RVT U4445 ( .A1(n4588), .A2(n276), .Y(n4583) );
  AND2X1_RVT U4446 ( .A1(n4377), .A2(n4254), .Y(n4588) );
  OR2X1_RVT U4447 ( .A1(n4103), .A2(n4589), .Y(n4254) );
  OR2X1_RVT U4448 ( .A1(n12722), .A2(n12512), .Y(n4589) );
  AND4X1_RVT U4449 ( .A1(n4271), .A2(n4590), .A3(n4463), .A4(n4591), .Y(n4554)
         );
  AND4X1_RVT U4450 ( .A1(n4592), .A2(n4593), .A3(n4594), .A4(n4595), .Y(n4591)
         );
  OR2X1_RVT U4451 ( .A1(n4234), .A2(n4155), .Y(n4595) );
  OR2X1_RVT U4452 ( .A1(n4172), .A2(n4201), .Y(n4594) );
  OR2X1_RVT U4453 ( .A1(n12710), .A2(n4426), .Y(n4593) );
  OR2X1_RVT U4454 ( .A1(n4150), .A2(n4132), .Y(n4426) );
  OR2X1_RVT U4455 ( .A1(n12718), .A2(n4214), .Y(n4132) );
  OR2X1_RVT U4456 ( .A1(n12526), .A2(n4255), .Y(n4592) );
  OR2X1_RVT U4457 ( .A1(n4136), .A2(n4364), .Y(n4255) );
  OR2X1_RVT U4458 ( .A1(n12510), .A2(n4340), .Y(n4364) );
  AND2X1_RVT U4459 ( .A1(n4596), .A2(n4597), .Y(n4463) );
  OR2X1_RVT U4460 ( .A1(n4598), .A2(n4203), .Y(n4597) );
  OR2X1_RVT U4461 ( .A1(n12536), .A2(n276), .Y(n4598) );
  OR2X1_RVT U4462 ( .A1(n4599), .A2(n4086), .Y(n4596) );
  OR2X1_RVT U4463 ( .A1(n12709), .A2(n4203), .Y(n4086) );
  OR2X1_RVT U4464 ( .A1(n4100), .A2(n4150), .Y(n4599) );
  OR2X1_RVT U4465 ( .A1(n12518), .A2(n4469), .Y(n4590) );
  AND2X1_RVT U4466 ( .A1(n4600), .A2(n4601), .Y(n4271) );
  OR2X1_RVT U4467 ( .A1(n4154), .A2(n4192), .Y(n4601) );
  OR2X1_RVT U4468 ( .A1(n4602), .A2(n4603), .Y(n4600) );
  AND4X1_RVT U4469 ( .A1(n4604), .A2(n4605), .A3(n4606), .A4(n4607), .Y(n4553)
         );
  OR2X1_RVT U4470 ( .A1(n4608), .A2(n4340), .Y(n4607) );
  AND2X1_RVT U4471 ( .A1(n4609), .A2(n4349), .Y(n4608) );
  OR2X1_RVT U4472 ( .A1(n12524), .A2(n4565), .Y(n4349) );
  OR2X1_RVT U4473 ( .A1(n4610), .A2(n12715), .Y(n4606) );
  AND2X1_RVT U4474 ( .A1(n4277), .A2(n4242), .Y(n4610) );
  OR2X1_RVT U4475 ( .A1(n12709), .A2(n4218), .Y(n4242) );
  OR2X1_RVT U4476 ( .A1(n4611), .A2(n4297), .Y(n4605) );
  AND2X1_RVT U4477 ( .A1(n4612), .A2(n4613), .Y(n4611) );
  OR2X1_RVT U4478 ( .A1(n12513), .A2(n4156), .Y(n4613) );
  AND2X1_RVT U4479 ( .A1(n4614), .A2(n4194), .Y(n4612) );
  OR2X1_RVT U4480 ( .A1(n274), .A2(n4153), .Y(n4614) );
  OR2X1_RVT U4481 ( .A1(n4615), .A2(n4094), .Y(n4604) );
  AND2X1_RVT U4482 ( .A1(n4616), .A2(n4617), .Y(n4615) );
  NAND2X1_RVT U4483 ( .A1(n4079), .A2(n4457), .Y(n4617) );
  AND2X1_RVT U4484 ( .A1(n4618), .A2(n4307), .Y(n4616) );
  OR2X1_RVT U4485 ( .A1(n4240), .A2(n4565), .Y(n4307) );
  OR2X1_RVT U4486 ( .A1(n12533), .A2(n4619), .Y(n4618) );
  AND4X1_RVT U4487 ( .A1(n4620), .A2(n4621), .A3(n4622), .A4(n4623), .Y(n4552)
         );
  OR2X1_RVT U4488 ( .A1(n4624), .A2(n4117), .Y(n4623) );
  AND2X1_RVT U4489 ( .A1(n4625), .A2(n4258), .Y(n4624) );
  AND2X1_RVT U4490 ( .A1(n4626), .A2(n4280), .Y(n4625) );
  OR2X1_RVT U4491 ( .A1(n276), .A2(n4603), .Y(n4280) );
  OR2X1_RVT U4492 ( .A1(n12512), .A2(n4214), .Y(n4603) );
  OR2X1_RVT U4493 ( .A1(n4627), .A2(n12529), .Y(n4622) );
  AND2X1_RVT U4494 ( .A1(n4628), .A2(n4629), .Y(n4627) );
  OR2X1_RVT U4495 ( .A1(n4630), .A2(n12707), .Y(n4629) );
  AND2X1_RVT U4496 ( .A1(n4631), .A2(n4632), .Y(n4630) );
  OR2X1_RVT U4497 ( .A1(n12511), .A2(n4491), .Y(n4632) );
  OR2X1_RVT U4498 ( .A1(n12714), .A2(n4137), .Y(n4631) );
  AND2X1_RVT U4499 ( .A1(n4633), .A2(n4634), .Y(n4628) );
  OR2X1_RVT U4500 ( .A1(n4103), .A2(n4635), .Y(n4633) );
  OR2X1_RVT U4501 ( .A1(n4636), .A2(n4137), .Y(n4621) );
  AND4X1_RVT U4502 ( .A1(n4637), .A2(n4638), .A3(n4639), .A4(n4103), .Y(n4636)
         );
  OR2X1_RVT U4503 ( .A1(n12715), .A2(n4153), .Y(n4639) );
  OR2X1_RVT U4504 ( .A1(n12523), .A2(n4172), .Y(n4638) );
  OR2X1_RVT U4505 ( .A1(n4225), .A2(n4203), .Y(n4637) );
  OR2X1_RVT U4506 ( .A1(n4640), .A2(n4079), .Y(n4620) );
  AND4X1_RVT U4507 ( .A1(n4504), .A2(n4641), .A3(n4302), .A4(n4218), .Y(n4640)
         );
  OR2X1_RVT U4508 ( .A1(n4172), .A2(n4635), .Y(n4302) );
  OR2X1_RVT U4509 ( .A1(n4340), .A2(n4547), .Y(n4641) );
  OR2X1_RVT U4510 ( .A1(n12517), .A2(n4305), .Y(n4504) );
  AND4X1_RVT U4511 ( .A1(n4643), .A2(n4644), .A3(n4645), .A4(n4646), .Y(n4642)
         );
  AND4X1_RVT U4512 ( .A1(n4155), .A2(n4391), .A3(n4647), .A4(n4648), .Y(n4646)
         );
  AND4X1_RVT U4513 ( .A1(n4470), .A2(n4415), .A3(n4560), .A4(n4561), .Y(n4648)
         );
  OR2X1_RVT U4514 ( .A1(n4563), .A2(n4076), .Y(n4561) );
  OR2X1_RVT U4515 ( .A1(n12713), .A2(n4194), .Y(n4076) );
  OR2X1_RVT U4516 ( .A1(n4093), .A2(n4602), .Y(n4560) );
  OR2X1_RVT U4517 ( .A1(n12718), .A2(n12531), .Y(n4602) );
  OR2X1_RVT U4518 ( .A1(n12707), .A2(n4214), .Y(n4093) );
  OR2X1_RVT U4519 ( .A1(n12719), .A2(n4112), .Y(n4415) );
  OR2X1_RVT U4520 ( .A1(n12540), .A2(n12524), .Y(n4112) );
  OR2X1_RVT U4521 ( .A1(n4234), .A2(n4649), .Y(n4470) );
  OR2X1_RVT U4522 ( .A1(n12531), .A2(n4138), .Y(n4649) );
  OR2X1_RVT U4523 ( .A1(n4136), .A2(n4650), .Y(n4647) );
  OR2X1_RVT U4524 ( .A1(n4264), .A2(n12522), .Y(n4650) );
  OR2X1_RVT U4525 ( .A1(n4203), .A2(n4651), .Y(n4391) );
  OR2X1_RVT U4526 ( .A1(n4137), .A2(n12529), .Y(n4651) );
  OR2X1_RVT U4527 ( .A1(n12711), .A2(n4562), .Y(n4155) );
  OR2X1_RVT U4528 ( .A1(n12524), .A2(n4154), .Y(n4562) );
  AND4X1_RVT U4529 ( .A1(n4652), .A2(n4653), .A3(n4654), .A4(n4655), .Y(n4645)
         );
  AND4X1_RVT U4530 ( .A1(n4656), .A2(n4657), .A3(n4658), .A4(n4659), .Y(n4655)
         );
  OR2X1_RVT U4531 ( .A1(n4170), .A2(n4660), .Y(n4659) );
  OR2X1_RVT U4532 ( .A1(n12513), .A2(n4240), .Y(n4660) );
  OR2X1_RVT U4533 ( .A1(n4153), .A2(n4661), .Y(n4658) );
  OR2X1_RVT U4534 ( .A1(n4662), .A2(n4117), .Y(n4661) );
  AND2X1_RVT U4535 ( .A1(n4096), .A2(n4156), .Y(n4662) );
  OR2X1_RVT U4536 ( .A1(n4663), .A2(n4664), .Y(n4657) );
  AND2X1_RVT U4537 ( .A1(n4311), .A2(n4267), .Y(n4663) );
  OR2X1_RVT U4538 ( .A1(n12712), .A2(n284), .Y(n4267) );
  OR2X1_RVT U4539 ( .A1(n12708), .A2(n12534), .Y(n4311) );
  OR2X1_RVT U4540 ( .A1(n4665), .A2(n4151), .Y(n4656) );
  AND2X1_RVT U4541 ( .A1(n4547), .A2(n4666), .Y(n4665) );
  OR2X1_RVT U4542 ( .A1(n12710), .A2(n276), .Y(n4666) );
  OR2X1_RVT U4543 ( .A1(n4667), .A2(n12536), .Y(n4654) );
  AND2X1_RVT U4544 ( .A1(n4538), .A2(n4668), .Y(n4667) );
  OR2X1_RVT U4545 ( .A1(n4144), .A2(n4491), .Y(n4668) );
  OR2X1_RVT U4546 ( .A1(n12517), .A2(n4356), .Y(n4538) );
  OR2X1_RVT U4547 ( .A1(n12714), .A2(n4144), .Y(n4356) );
  OR2X1_RVT U4548 ( .A1(n4669), .A2(n4305), .Y(n4653) );
  AND2X1_RVT U4549 ( .A1(n4258), .A2(n4530), .Y(n4669) );
  OR2X1_RVT U4550 ( .A1(n4114), .A2(n4203), .Y(n4258) );
  OR2X1_RVT U4551 ( .A1(n4670), .A2(n4194), .Y(n4652) );
  AND2X1_RVT U4552 ( .A1(n4157), .A2(n4159), .Y(n4670) );
  AND4X1_RVT U4553 ( .A1(n4671), .A2(n4672), .A3(n4673), .A4(n4674), .Y(n4644)
         );
  AND4X1_RVT U4554 ( .A1(n4675), .A2(n4676), .A3(n4677), .A4(n4678), .Y(n4674)
         );
  OR2X1_RVT U4555 ( .A1(n4679), .A2(n12520), .Y(n4678) );
  AND2X1_RVT U4556 ( .A1(n4085), .A2(n4377), .Y(n4679) );
  OR2X1_RVT U4557 ( .A1(n4234), .A2(n4265), .Y(n4377) );
  OR2X1_RVT U4558 ( .A1(n12523), .A2(n4117), .Y(n4265) );
  OR2X1_RVT U4559 ( .A1(n12527), .A2(n4680), .Y(n4085) );
  OR2X1_RVT U4560 ( .A1(n12510), .A2(n12516), .Y(n4680) );
  OR2X1_RVT U4561 ( .A1(n4681), .A2(n12534), .Y(n4677) );
  AND2X1_RVT U4562 ( .A1(n4394), .A2(n4682), .Y(n4681) );
  OR2X1_RVT U4563 ( .A1(n12539), .A2(n274), .Y(n4682) );
  OR2X1_RVT U4564 ( .A1(n12537), .A2(n4201), .Y(n4394) );
  OR2X1_RVT U4565 ( .A1(n4683), .A2(n12515), .Y(n4676) );
  AND2X1_RVT U4566 ( .A1(n4412), .A2(n4684), .Y(n4683) );
  OR2X1_RVT U4567 ( .A1(n12540), .A2(n4137), .Y(n4684) );
  OR2X1_RVT U4568 ( .A1(n4079), .A2(n4685), .Y(n4412) );
  OR2X1_RVT U4569 ( .A1(n4686), .A2(n4138), .Y(n4675) );
  AND2X1_RVT U4570 ( .A1(n4687), .A2(n4688), .Y(n4686) );
  OR2X1_RVT U4571 ( .A1(n4194), .A2(n12537), .Y(n4688) );
  AND2X1_RVT U4572 ( .A1(n4689), .A2(n4170), .Y(n4687) );
  OR2X1_RVT U4573 ( .A1(n4156), .A2(n4117), .Y(n4170) );
  OR2X1_RVT U4574 ( .A1(n12512), .A2(n4201), .Y(n4689) );
  OR2X1_RVT U4575 ( .A1(n12722), .A2(n4156), .Y(n4201) );
  OR2X1_RVT U4576 ( .A1(n4690), .A2(n4214), .Y(n4673) );
  AND4X1_RVT U4577 ( .A1(n4691), .A2(n4692), .A3(n4367), .A4(n4277), .Y(n4690)
         );
  OR2X1_RVT U4578 ( .A1(n4340), .A2(n4440), .Y(n4277) );
  OR2X1_RVT U4579 ( .A1(n4172), .A2(n4619), .Y(n4367) );
  OR2X1_RVT U4580 ( .A1(n12518), .A2(n12511), .Y(n4619) );
  OR2X1_RVT U4581 ( .A1(n276), .A2(n4094), .Y(n4692) );
  OR2X1_RVT U4582 ( .A1(n274), .A2(n12537), .Y(n4691) );
  OR2X1_RVT U4583 ( .A1(n4693), .A2(n4150), .Y(n4672) );
  AND2X1_RVT U4584 ( .A1(n4694), .A2(n4171), .Y(n4693) );
  AND2X1_RVT U4585 ( .A1(n4626), .A2(n4421), .Y(n4694) );
  OR2X1_RVT U4586 ( .A1(n4695), .A2(n12719), .Y(n4421) );
  AND2X1_RVT U4587 ( .A1(n4192), .A2(n4696), .Y(n4695) );
  OR2X1_RVT U4588 ( .A1(n12515), .A2(n4079), .Y(n4696) );
  OR2X1_RVT U4589 ( .A1(n4240), .A2(n4378), .Y(n4626) );
  OR2X1_RVT U4590 ( .A1(n4225), .A2(n4114), .Y(n4378) );
  OR2X1_RVT U4591 ( .A1(n4697), .A2(n4218), .Y(n4671) );
  AND2X1_RVT U4592 ( .A1(n4698), .A2(n12523), .Y(n4697) );
  AND2X1_RVT U4593 ( .A1(n4699), .A2(n4399), .Y(n4698) );
  OR2X1_RVT U4594 ( .A1(n4240), .A2(n4340), .Y(n4699) );
  AND4X1_RVT U4595 ( .A1(n4700), .A2(n4701), .A3(n4702), .A4(n4703), .Y(n4643)
         );
  AND2X1_RVT U4596 ( .A1(n4704), .A2(n4705), .Y(n4703) );
  OR2X1_RVT U4597 ( .A1(n12715), .A2(n4320), .Y(n4705) );
  OR2X1_RVT U4598 ( .A1(n12531), .A2(n4706), .Y(n4320) );
  OR2X1_RVT U4599 ( .A1(n4136), .A2(n4225), .Y(n4706) );
  AND2X1_RVT U4600 ( .A1(n4707), .A2(n4708), .Y(n4704) );
  OR2X1_RVT U4601 ( .A1(n4109), .A2(n4120), .Y(n4708) );
  OR2X1_RVT U4602 ( .A1(n4153), .A2(n4348), .Y(n4120) );
  OR2X1_RVT U4603 ( .A1(n12711), .A2(n4114), .Y(n4348) );
  OR2X1_RVT U4604 ( .A1(n4156), .A2(n4233), .Y(n4707) );
  OR2X1_RVT U4605 ( .A1(n4144), .A2(n4709), .Y(n4233) );
  OR2X1_RVT U4606 ( .A1(n4144), .A2(n4324), .Y(n4702) );
  OR2X1_RVT U4607 ( .A1(n276), .A2(n12533), .Y(n4324) );
  OR2X1_RVT U4608 ( .A1(n4710), .A2(n4100), .Y(n4701) );
  AND4X1_RVT U4609 ( .A1(n4711), .A2(n4712), .A3(n4713), .A4(n4714), .Y(n4710)
         );
  OR2X1_RVT U4610 ( .A1(n12709), .A2(n4715), .Y(n4713) );
  OR2X1_RVT U4611 ( .A1(n4716), .A2(n12716), .Y(n4715) );
  AND2X1_RVT U4612 ( .A1(n4151), .A2(n4717), .Y(n4716) );
  OR2X1_RVT U4613 ( .A1(n12526), .A2(n4718), .Y(n4712) );
  OR2X1_RVT U4614 ( .A1(n4457), .A2(n4094), .Y(n4718) );
  OR2X1_RVT U4615 ( .A1(n4077), .A2(n4103), .Y(n4711) );
  OR2X1_RVT U4616 ( .A1(n12713), .A2(n4203), .Y(n4103) );
  OR2X1_RVT U4617 ( .A1(n4577), .A2(n4491), .Y(n4700) );
  OR2X1_RVT U4618 ( .A1(n12542), .A2(n4114), .Y(n4491) );
  AND4X1_RVT U4619 ( .A1(n4720), .A2(n4721), .A3(n4722), .A4(n4723), .Y(n4719)
         );
  AND4X1_RVT U4620 ( .A1(n4724), .A2(n4725), .A3(n4726), .A4(n4727), .Y(n4723)
         );
  AND4X1_RVT U4621 ( .A1(n4728), .A2(n4729), .A3(n4730), .A4(n4731), .Y(n4727)
         );
  OR2X1_RVT U4622 ( .A1(n4565), .A2(n4709), .Y(n4731) );
  OR2X1_RVT U4623 ( .A1(n12712), .A2(n12536), .Y(n4709) );
  OR2X1_RVT U4624 ( .A1(n12510), .A2(n12520), .Y(n4565) );
  OR2X1_RVT U4625 ( .A1(n4732), .A2(n4151), .Y(n4730) );
  AND2X1_RVT U4626 ( .A1(n4097), .A2(n4664), .Y(n4732) );
  OR2X1_RVT U4627 ( .A1(n276), .A2(n4733), .Y(n4097) );
  OR2X1_RVT U4628 ( .A1(n12510), .A2(n12709), .Y(n4733) );
  OR2X1_RVT U4629 ( .A1(n4734), .A2(n4079), .Y(n4729) );
  OR2X1_RVT U4630 ( .A1(n12524), .A2(n4240), .Y(n4079) );
  AND2X1_RVT U4631 ( .A1(n4215), .A2(n4735), .Y(n4734) );
  OR2X1_RVT U4632 ( .A1(n4094), .A2(n4296), .Y(n4735) );
  OR2X1_RVT U4633 ( .A1(n12528), .A2(n12516), .Y(n4094) );
  OR2X1_RVT U4634 ( .A1(n4340), .A2(n4736), .Y(n4215) );
  OR2X1_RVT U4635 ( .A1(n12720), .A2(n12531), .Y(n4736) );
  OR2X1_RVT U4636 ( .A1(n4737), .A2(n4138), .Y(n4728) );
  AND2X1_RVT U4637 ( .A1(n4535), .A2(n4738), .Y(n4737) );
  OR2X1_RVT U4638 ( .A1(n4739), .A2(n12709), .Y(n4738) );
  AND2X1_RVT U4639 ( .A1(n4194), .A2(n4547), .Y(n4739) );
  OR2X1_RVT U4640 ( .A1(n12717), .A2(n4156), .Y(n4547) );
  OR2X1_RVT U4641 ( .A1(n12537), .A2(n4740), .Y(n4535) );
  OR2X1_RVT U4642 ( .A1(n12722), .A2(n12718), .Y(n4740) );
  OR2X1_RVT U4643 ( .A1(n4741), .A2(n12515), .Y(n4726) );
  AND2X1_RVT U4644 ( .A1(n4742), .A2(n4743), .Y(n4741) );
  OR2X1_RVT U4645 ( .A1(n4744), .A2(n4240), .Y(n4743) );
  AND2X1_RVT U4646 ( .A1(n4305), .A2(n4745), .Y(n4744) );
  OR2X1_RVT U4647 ( .A1(n4096), .A2(n4218), .Y(n4742) );
  OR2X1_RVT U4648 ( .A1(n12529), .A2(n4154), .Y(n4218) );
  OR2X1_RVT U4649 ( .A1(n4746), .A2(n12718), .Y(n4725) );
  AND2X1_RVT U4650 ( .A1(n4310), .A2(n4469), .Y(n4746) );
  OR2X1_RVT U4651 ( .A1(n12527), .A2(n4747), .Y(n4469) );
  OR2X1_RVT U4652 ( .A1(n4150), .A2(n12516), .Y(n4747) );
  OR2X1_RVT U4653 ( .A1(n4096), .A2(n4577), .Y(n4310) );
  OR2X1_RVT U4654 ( .A1(n12516), .A2(n12531), .Y(n4577) );
  OR2X1_RVT U4655 ( .A1(n4748), .A2(n12513), .Y(n4724) );
  AND2X1_RVT U4656 ( .A1(n4350), .A2(n4749), .Y(n4748) );
  OR2X1_RVT U4657 ( .A1(n4564), .A2(n4144), .Y(n4749) );
  OR2X1_RVT U4658 ( .A1(n4203), .A2(n4685), .Y(n4350) );
  OR2X1_RVT U4659 ( .A1(n12717), .A2(n276), .Y(n4685) );
  AND2X1_RVT U4660 ( .A1(n12517), .A2(n12720), .Y(n4446) );
  AND4X1_RVT U4661 ( .A1(n4750), .A2(n4751), .A3(n4752), .A4(n4753), .Y(n4722)
         );
  AND4X1_RVT U4662 ( .A1(n4754), .A2(n4755), .A3(n4756), .A4(n4757), .Y(n4753)
         );
  OR2X1_RVT U4663 ( .A1(n4758), .A2(n12522), .Y(n4757) );
  AND2X1_RVT U4664 ( .A1(n4337), .A2(n4408), .Y(n4758) );
  OR2X1_RVT U4665 ( .A1(n4153), .A2(n4664), .Y(n4408) );
  OR2X1_RVT U4666 ( .A1(n12720), .A2(n4150), .Y(n4664) );
  OR2X1_RVT U4667 ( .A1(n12707), .A2(n12512), .Y(n4153) );
  OR2X1_RVT U4668 ( .A1(n12513), .A2(n4440), .Y(n4337) );
  OR2X1_RVT U4669 ( .A1(n12517), .A2(n12531), .Y(n4440) );
  OR2X1_RVT U4670 ( .A1(n4759), .A2(n12716), .Y(n4756) );
  AND2X1_RVT U4671 ( .A1(n4499), .A2(n4760), .Y(n4759) );
  OR2X1_RVT U4672 ( .A1(n4457), .A2(n4167), .Y(n4760) );
  OR2X1_RVT U4673 ( .A1(n4340), .A2(n4761), .Y(n4167) );
  OR2X1_RVT U4674 ( .A1(n12542), .A2(n12518), .Y(n4761) );
  OR2X1_RVT U4675 ( .A1(n12526), .A2(n4762), .Y(n4499) );
  OR2X1_RVT U4676 ( .A1(n4340), .A2(n4136), .Y(n4762) );
  OR2X1_RVT U4677 ( .A1(n4763), .A2(n12722), .Y(n4755) );
  AND2X1_RVT U4678 ( .A1(n4445), .A2(n4374), .Y(n4763) );
  OR2X1_RVT U4679 ( .A1(n4156), .A2(n4192), .Y(n4374) );
  OR2X1_RVT U4680 ( .A1(n12714), .A2(n4340), .Y(n4192) );
  OR2X1_RVT U4681 ( .A1(n4564), .A2(n4172), .Y(n4445) );
  OR2X1_RVT U4682 ( .A1(n12523), .A2(n12719), .Y(n4564) );
  OR2X1_RVT U4683 ( .A1(n4764), .A2(n4214), .Y(n4754) );
  AND2X1_RVT U4684 ( .A1(n4765), .A2(n4766), .Y(n4764) );
  OR2X1_RVT U4685 ( .A1(n4136), .A2(n4563), .Y(n4766) );
  OR2X1_RVT U4686 ( .A1(n12716), .A2(n284), .Y(n4563) );
  AND2X1_RVT U4687 ( .A1(n4767), .A2(n4431), .Y(n4765) );
  OR2X1_RVT U4688 ( .A1(n4144), .A2(n4768), .Y(n4431) );
  OR2X1_RVT U4689 ( .A1(n12539), .A2(n12518), .Y(n4768) );
  OR2X1_RVT U4690 ( .A1(n4200), .A2(n4137), .Y(n4752) );
  OR2X1_RVT U4691 ( .A1(n12709), .A2(n4096), .Y(n4200) );
  OR2X1_RVT U4692 ( .A1(n4769), .A2(n4100), .Y(n4751) );
  AND2X1_RVT U4693 ( .A1(n4770), .A2(n4281), .Y(n4769) );
  AND2X1_RVT U4694 ( .A1(n4771), .A2(n4772), .Y(n4281) );
  OR2X1_RVT U4695 ( .A1(n12527), .A2(n4305), .Y(n4772) );
  OR2X1_RVT U4696 ( .A1(n4203), .A2(n4077), .Y(n4771) );
  OR2X1_RVT U4697 ( .A1(n12512), .A2(n4150), .Y(n4077) );
  AND2X1_RVT U4698 ( .A1(n4773), .A2(n4467), .Y(n4770) );
  OR2X1_RVT U4699 ( .A1(n4234), .A2(n4717), .Y(n4467) );
  OR2X1_RVT U4700 ( .A1(n12711), .A2(n274), .Y(n4717) );
  OR2X1_RVT U4701 ( .A1(n4096), .A2(n4263), .Y(n4773) );
  OR2X1_RVT U4702 ( .A1(n12511), .A2(n4774), .Y(n4263) );
  OR2X1_RVT U4703 ( .A1(n12707), .A2(n12540), .Y(n4774) );
  OR2X1_RVT U4704 ( .A1(n4775), .A2(n12707), .Y(n4750) );
  AND4X1_RVT U4705 ( .A1(n4776), .A2(n4777), .A3(n4778), .A4(n4609), .Y(n4775)
         );
  OR2X1_RVT U4706 ( .A1(n4150), .A2(n4530), .Y(n4609) );
  OR2X1_RVT U4707 ( .A1(n12712), .A2(n12718), .Y(n4530) );
  OR2X1_RVT U4708 ( .A1(n4150), .A2(n4779), .Y(n4778) );
  OR2X1_RVT U4709 ( .A1(n12517), .A2(n12522), .Y(n4779) );
  OR2X1_RVT U4710 ( .A1(n12717), .A2(n4109), .Y(n4150) );
  OR2X1_RVT U4711 ( .A1(n4780), .A2(n4231), .Y(n4777) );
  OR2X1_RVT U4712 ( .A1(n12511), .A2(n4075), .Y(n4231) );
  AND2X1_RVT U4713 ( .A1(n4214), .A2(n4781), .Y(n4780) );
  OR2X1_RVT U4714 ( .A1(n12715), .A2(n4114), .Y(n4781) );
  OR2X1_RVT U4715 ( .A1(n12711), .A2(n12522), .Y(n4214) );
  OR2X1_RVT U4716 ( .A1(n12713), .A2(n4745), .Y(n4776) );
  OR2X1_RVT U4717 ( .A1(n12717), .A2(n4154), .Y(n4745) );
  OR2X1_RVT U4718 ( .A1(n4100), .A2(n274), .Y(n4154) );
  AND4X1_RVT U4719 ( .A1(n4782), .A2(n4783), .A3(n4784), .A4(n4785), .Y(n4721)
         );
  AND4X1_RVT U4720 ( .A1(n4786), .A2(n4787), .A3(n4788), .A4(n4789), .Y(n4785)
         );
  OR2X1_RVT U4721 ( .A1(n4172), .A2(n4299), .Y(n4789) );
  OR2X1_RVT U4722 ( .A1(n12524), .A2(n4194), .Y(n4299) );
  OR2X1_RVT U4723 ( .A1(n12528), .A2(n4340), .Y(n4172) );
  OR2X1_RVT U4724 ( .A1(n4159), .A2(n4635), .Y(n4788) );
  OR2X1_RVT U4725 ( .A1(n12721), .A2(n12511), .Y(n4635) );
  OR2X1_RVT U4726 ( .A1(n4225), .A2(n4151), .Y(n4159) );
  OR2X1_RVT U4727 ( .A1(n4144), .A2(n4171), .Y(n4787) );
  OR2X1_RVT U4728 ( .A1(n12520), .A2(n12533), .Y(n4171) );
  OR2X1_RVT U4729 ( .A1(n12510), .A2(n12708), .Y(n4144) );
  OR2X1_RVT U4730 ( .A1(n284), .A2(n4510), .Y(n4786) );
  OR2X1_RVT U4731 ( .A1(n12518), .A2(n4297), .Y(n4510) );
  OR2X1_RVT U4732 ( .A1(n4114), .A2(n4544), .Y(n4784) );
  OR2X1_RVT U4733 ( .A1(n284), .A2(n4790), .Y(n4544) );
  OR2X1_RVT U4734 ( .A1(n12714), .A2(n12531), .Y(n4790) );
  AND2X1_RVT U4735 ( .A1(n12512), .A2(n12515), .Y(n4574) );
  OR2X1_RVT U4736 ( .A1(n4156), .A2(n4104), .Y(n4783) );
  OR2X1_RVT U4737 ( .A1(n12540), .A2(n4791), .Y(n4104) );
  OR2X1_RVT U4738 ( .A1(n12715), .A2(n12707), .Y(n4791) );
  OR2X1_RVT U4739 ( .A1(n12517), .A2(n4136), .Y(n4156) );
  OR2X1_RVT U4740 ( .A1(n4203), .A2(n4767), .Y(n4782) );
  OR2X1_RVT U4741 ( .A1(n12513), .A2(n4158), .Y(n4767) );
  OR2X1_RVT U4742 ( .A1(n12717), .A2(n12718), .Y(n4158) );
  AND4X1_RVT U4743 ( .A1(n4792), .A2(n4269), .A3(n4793), .A4(n4794), .Y(n4720)
         );
  OR2X1_RVT U4744 ( .A1(n12517), .A2(n4714), .Y(n4794) );
  OR2X1_RVT U4745 ( .A1(n12713), .A2(n4264), .Y(n4714) );
  OR2X1_RVT U4746 ( .A1(n12515), .A2(n4305), .Y(n4264) );
  OR2X1_RVT U4747 ( .A1(n12510), .A2(n4131), .Y(n4305) );
  AND2X1_RVT U4748 ( .A1(n4795), .A2(n4796), .Y(n4793) );
  OR2X1_RVT U4749 ( .A1(n12539), .A2(n4634), .Y(n4796) );
  OR2X1_RVT U4750 ( .A1(n4203), .A2(n4296), .Y(n4634) );
  OR2X1_RVT U4751 ( .A1(n12517), .A2(n12511), .Y(n4296) );
  OR2X1_RVT U4752 ( .A1(n12512), .A2(n4092), .Y(n4131) );
  OR2X1_RVT U4753 ( .A1(n12720), .A2(n4365), .Y(n4795) );
  OR2X1_RVT U4754 ( .A1(n12536), .A2(n4399), .Y(n4365) );
  OR2X1_RVT U4755 ( .A1(n12712), .A2(n12707), .Y(n4399) );
  OR2X1_RVT U4756 ( .A1(n12710), .A2(n12528), .Y(n4075) );
  AND2X1_RVT U4757 ( .A1(n4797), .A2(n4798), .Y(n4269) );
  OR2X1_RVT U4758 ( .A1(n4151), .A2(n4137), .Y(n4798) );
  OR2X1_RVT U4759 ( .A1(n12719), .A2(n4109), .Y(n4137) );
  AND2X1_RVT U4760 ( .A1(n4136), .A2(n4100), .Y(n4189) );
  OR2X1_RVT U4761 ( .A1(n12523), .A2(n4203), .Y(n4151) );
  OR2X1_RVT U4762 ( .A1(n12708), .A2(n4240), .Y(n4203) );
  OR2X1_RVT U4763 ( .A1(n4799), .A2(n4194), .Y(n4797) );
  OR2X1_RVT U4764 ( .A1(n12517), .A2(n274), .Y(n4194) );
  AND2X1_RVT U4765 ( .A1(n12721), .A2(n12510), .Y(n4457) );
  OR2X1_RVT U4766 ( .A1(n12516), .A2(n4297), .Y(n4799) );
  OR2X1_RVT U4767 ( .A1(n12717), .A2(n12533), .Y(n4297) );
  AND2X1_RVT U4768 ( .A1(n4800), .A2(n4801), .Y(n4792) );
  OR2X1_RVT U4769 ( .A1(n4117), .A2(n4450), .Y(n4801) );
  OR2X1_RVT U4770 ( .A1(n12518), .A2(n4157), .Y(n4450) );
  OR2X1_RVT U4771 ( .A1(n12533), .A2(n4234), .Y(n4157) );
  OR2X1_RVT U4772 ( .A1(n12513), .A2(n12516), .Y(n4234) );
  OR2X1_RVT U4773 ( .A1(n12714), .A2(n12712), .Y(n4096) );
  OR2X1_RVT U4774 ( .A1(n12722), .A2(n12716), .Y(n4117) );
  XOR2X1_RVT U4775 ( .A1(key[20]), .A2(state[20]), .Y(n4092) );
  OR2X1_RVT U4776 ( .A1(n4109), .A2(n4238), .Y(n4800) );
  OR2X1_RVT U4777 ( .A1(n4340), .A2(n4531), .Y(n4238) );
  OR2X1_RVT U4778 ( .A1(n12520), .A2(n4138), .Y(n4531) );
  OR2X1_RVT U4779 ( .A1(n12715), .A2(n4240), .Y(n4138) );
  XOR2X1_RVT U4780 ( .A1(key[18]), .A2(state[18]), .Y(n4240) );
  XOR2X1_RVT U4781 ( .A1(key[19]), .A2(state[19]), .Y(n4174) );
  OR2X1_RVT U4782 ( .A1(n12720), .A2(n12518), .Y(n4114) );
  XOR2X1_RVT U4783 ( .A1(key[21]), .A2(state[21]), .Y(n4100) );
  XOR2X1_RVT U4784 ( .A1(key[22]), .A2(state[22]), .Y(n4136) );
  OR2X1_RVT U4785 ( .A1(n12710), .A2(n12516), .Y(n4340) );
  XOR2X1_RVT U4786 ( .A1(key[16]), .A2(state[16]), .Y(n4115) );
  XOR2X1_RVT U4787 ( .A1(key[17]), .A2(state[17]), .Y(n4225) );
  XOR2X1_RVT U4788 ( .A1(key[23]), .A2(state[23]), .Y(n4109) );
  AND4X1_RVT U4789 ( .A1(n4803), .A2(n4804), .A3(n4805), .A4(n4806), .Y(n4802)
         );
  AND4X1_RVT U4790 ( .A1(n4807), .A2(n4808), .A3(n4809), .A4(n4810), .Y(n4806)
         );
  AND4X1_RVT U4791 ( .A1(n4811), .A2(n4812), .A3(n4813), .A4(n4814), .Y(n4810)
         );
  OR2X1_RVT U4792 ( .A1(n12471), .A2(n4816), .Y(n4809) );
  OR2X1_RVT U4793 ( .A1(n4817), .A2(n4818), .Y(n4807) );
  OR2X1_RVT U4794 ( .A1(n12704), .A2(n4819), .Y(n4818) );
  AND4X1_RVT U4795 ( .A1(n4820), .A2(n4821), .A3(n4822), .A4(n4823), .Y(n4805)
         );
  OR2X1_RVT U4796 ( .A1(n4824), .A2(n12702), .Y(n4823) );
  AND2X1_RVT U4797 ( .A1(n4825), .A2(n4826), .Y(n4824) );
  AND2X1_RVT U4798 ( .A1(n4827), .A2(n4828), .Y(n4822) );
  OR2X1_RVT U4799 ( .A1(n4829), .A2(n296), .Y(n4828) );
  AND2X1_RVT U4800 ( .A1(n4830), .A2(n4831), .Y(n4829) );
  OR2X1_RVT U4801 ( .A1(n12462), .A2(n4833), .Y(n4831) );
  OR2X1_RVT U4802 ( .A1(n4819), .A2(n4834), .Y(n4830) );
  OR2X1_RVT U4803 ( .A1(n4835), .A2(n12468), .Y(n4827) );
  AND2X1_RVT U4804 ( .A1(n4837), .A2(n4838), .Y(n4835) );
  OR2X1_RVT U4805 ( .A1(n4839), .A2(n4840), .Y(n4821) );
  AND2X1_RVT U4806 ( .A1(n4841), .A2(n4842), .Y(n4839) );
  OR2X1_RVT U4807 ( .A1(n12463), .A2(n4843), .Y(n4842) );
  AND2X1_RVT U4808 ( .A1(n4844), .A2(n4845), .Y(n4841) );
  AND2X1_RVT U4809 ( .A1(n4846), .A2(n4847), .Y(n4820) );
  OR2X1_RVT U4810 ( .A1(n4848), .A2(n12445), .Y(n4847) );
  AND2X1_RVT U4811 ( .A1(n4850), .A2(n4851), .Y(n4848) );
  OR2X1_RVT U4812 ( .A1(n4852), .A2(n4853), .Y(n4851) );
  OR2X1_RVT U4813 ( .A1(n12454), .A2(n12449), .Y(n4853) );
  OR2X1_RVT U4814 ( .A1(n4856), .A2(n4857), .Y(n4846) );
  AND2X1_RVT U4815 ( .A1(n4858), .A2(n4859), .Y(n4856) );
  AND2X1_RVT U4816 ( .A1(n4860), .A2(n4861), .Y(n4858) );
  AND4X1_RVT U4817 ( .A1(n4862), .A2(n4863), .A3(n4864), .A4(n4865), .Y(n4804)
         );
  AND4X1_RVT U4818 ( .A1(n4866), .A2(n4867), .A3(n4868), .A4(n4869), .Y(n4865)
         );
  OR2X1_RVT U4819 ( .A1(n4870), .A2(n12474), .Y(n4869) );
  AND4X1_RVT U4820 ( .A1(n4872), .A2(n4873), .A3(n4874), .A4(n4875), .Y(n4870)
         );
  OR2X1_RVT U4821 ( .A1(n4876), .A2(n4843), .Y(n4875) );
  OR2X1_RVT U4822 ( .A1(n4877), .A2(n12460), .Y(n4874) );
  OR2X1_RVT U4823 ( .A1(n4879), .A2(n12451), .Y(n4868) );
  AND4X1_RVT U4824 ( .A1(n4880), .A2(n4881), .A3(n4882), .A4(n4883), .Y(n4879)
         );
  OR2X1_RVT U4825 ( .A1(n4884), .A2(n4885), .Y(n4883) );
  OR2X1_RVT U4826 ( .A1(n12468), .A2(n12463), .Y(n4885) );
  AND2X1_RVT U4827 ( .A1(n4886), .A2(n4887), .Y(n4882) );
  OR2X1_RVT U4828 ( .A1(n12706), .A2(n4888), .Y(n4881) );
  OR2X1_RVT U4829 ( .A1(n4889), .A2(n4890), .Y(n4880) );
  AND2X1_RVT U4830 ( .A1(n4891), .A2(n4892), .Y(n4889) );
  OR2X1_RVT U4831 ( .A1(n12468), .A2(n4893), .Y(n4892) );
  OR2X1_RVT U4832 ( .A1(n4826), .A2(n4894), .Y(n4867) );
  OR2X1_RVT U4833 ( .A1(n4893), .A2(n4895), .Y(n4866) );
  OR2X1_RVT U4834 ( .A1(n4896), .A2(n4897), .Y(n4864) );
  OR2X1_RVT U4835 ( .A1(n4898), .A2(n4891), .Y(n4863) );
  OR2X1_RVT U4836 ( .A1(n4899), .A2(n4900), .Y(n4862) );
  AND4X1_RVT U4837 ( .A1(n4901), .A2(n4902), .A3(n4903), .A4(n4904), .Y(n4803)
         );
  AND2X1_RVT U4838 ( .A1(n4905), .A2(n4906), .Y(n4904) );
  OR2X1_RVT U4839 ( .A1(n4890), .A2(n4907), .Y(n4906) );
  AND2X1_RVT U4840 ( .A1(n4908), .A2(n4909), .Y(n4905) );
  OR2X1_RVT U4841 ( .A1(n4910), .A2(n4833), .Y(n4909) );
  OR2X1_RVT U4842 ( .A1(n4834), .A2(n4911), .Y(n4908) );
  OR2X1_RVT U4843 ( .A1(n294), .A2(n4912), .Y(n4903) );
  OR2X1_RVT U4844 ( .A1(n4913), .A2(n12458), .Y(n4902) );
  OR2X1_RVT U4845 ( .A1(n12461), .A2(n4915), .Y(n4901) );
  AND4X1_RVT U4846 ( .A1(n4917), .A2(n4918), .A3(n4919), .A4(n4920), .Y(n4916)
         );
  AND4X1_RVT U4847 ( .A1(n4921), .A2(n4812), .A3(n4922), .A4(n4923), .Y(n4920)
         );
  AND4X1_RVT U4848 ( .A1(n4924), .A2(n4925), .A3(n4926), .A4(n4927), .Y(n4923)
         );
  OR2X1_RVT U4849 ( .A1(n4833), .A2(n4928), .Y(n4927) );
  OR2X1_RVT U4850 ( .A1(n4929), .A2(n12473), .Y(n4928) );
  OR2X1_RVT U4851 ( .A1(n4834), .A2(n4930), .Y(n4926) );
  OR2X1_RVT U4852 ( .A1(n294), .A2(n12457), .Y(n4930) );
  OR2X1_RVT U4853 ( .A1(n4931), .A2(n4877), .Y(n4925) );
  AND2X1_RVT U4854 ( .A1(n4888), .A2(n4932), .Y(n4931) );
  OR2X1_RVT U4855 ( .A1(n4933), .A2(n4934), .Y(n4924) );
  AND2X1_RVT U4856 ( .A1(n4935), .A2(n4936), .Y(n4933) );
  AND2X1_RVT U4857 ( .A1(n4937), .A2(n4938), .Y(n4922) );
  OR2X1_RVT U4858 ( .A1(n4884), .A2(n4939), .Y(n4938) );
  OR2X1_RVT U4859 ( .A1(n4940), .A2(n12704), .Y(n4939) );
  OR2X1_RVT U4860 ( .A1(n4941), .A2(n4942), .Y(n4937) );
  OR2X1_RVT U4861 ( .A1(n4943), .A2(n12462), .Y(n4942) );
  OR2X1_RVT U4862 ( .A1(n4819), .A2(n4944), .Y(n4812) );
  AND4X1_RVT U4863 ( .A1(n4945), .A2(n4946), .A3(n4947), .A4(n4948), .Y(n4919)
         );
  AND4X1_RVT U4864 ( .A1(n4949), .A2(n4950), .A3(n4951), .A4(n4952), .Y(n4948)
         );
  OR2X1_RVT U4865 ( .A1(n4953), .A2(n12476), .Y(n4952) );
  AND2X1_RVT U4866 ( .A1(n4955), .A2(n4956), .Y(n4953) );
  OR2X1_RVT U4867 ( .A1(n12445), .A2(n4834), .Y(n4956) );
  OR2X1_RVT U4868 ( .A1(n4957), .A2(n4836), .Y(n4951) );
  AND2X1_RVT U4869 ( .A1(n4958), .A2(n4959), .Y(n4957) );
  OR2X1_RVT U4870 ( .A1(n4960), .A2(n12703), .Y(n4950) );
  AND2X1_RVT U4871 ( .A1(n4961), .A2(n4962), .Y(n4960) );
  OR2X1_RVT U4872 ( .A1(n4963), .A2(n4912), .Y(n4962) );
  AND2X1_RVT U4873 ( .A1(n12476), .A2(n12460), .Y(n4963) );
  OR2X1_RVT U4874 ( .A1(n4964), .A2(n12446), .Y(n4949) );
  AND2X1_RVT U4875 ( .A1(n4966), .A2(n4967), .Y(n4964) );
  OR2X1_RVT U4876 ( .A1(n4968), .A2(n12452), .Y(n4947) );
  AND2X1_RVT U4877 ( .A1(n4969), .A2(n4970), .Y(n4968) );
  OR2X1_RVT U4878 ( .A1(n12460), .A2(n4971), .Y(n4970) );
  AND2X1_RVT U4879 ( .A1(n4972), .A2(n4973), .Y(n4969) );
  OR2X1_RVT U4880 ( .A1(n4974), .A2(n4975), .Y(n4972) );
  OR2X1_RVT U4881 ( .A1(n4819), .A2(n4890), .Y(n4975) );
  OR2X1_RVT U4882 ( .A1(n4976), .A2(n12700), .Y(n4946) );
  AND2X1_RVT U4883 ( .A1(n4977), .A2(n4978), .Y(n4976) );
  OR2X1_RVT U4884 ( .A1(n4979), .A2(n4980), .Y(n4945) );
  AND2X1_RVT U4885 ( .A1(n4981), .A2(n4982), .Y(n4979) );
  AND2X1_RVT U4886 ( .A1(n4983), .A2(n4984), .Y(n4981) );
  OR2X1_RVT U4887 ( .A1(n296), .A2(n4912), .Y(n4984) );
  OR2X1_RVT U4888 ( .A1(n12470), .A2(n4877), .Y(n4983) );
  AND4X1_RVT U4889 ( .A1(n4985), .A2(n4986), .A3(n4987), .A4(n4988), .Y(n4918)
         );
  AND4X1_RVT U4890 ( .A1(n4989), .A2(n4990), .A3(n4991), .A4(n4992), .Y(n4988)
         );
  OR2X1_RVT U4891 ( .A1(n4912), .A2(n4911), .Y(n4992) );
  OR2X1_RVT U4892 ( .A1(n4843), .A2(n4993), .Y(n4991) );
  OR2X1_RVT U4893 ( .A1(n4876), .A2(n4994), .Y(n4990) );
  OR2X1_RVT U4894 ( .A1(n4819), .A2(n4995), .Y(n4989) );
  AND2X1_RVT U4895 ( .A1(n4996), .A2(n4997), .Y(n4987) );
  OR2X1_RVT U4896 ( .A1(n12471), .A2(n4998), .Y(n4997) );
  OR2X1_RVT U4897 ( .A1(n12450), .A2(n4895), .Y(n4996) );
  OR2X1_RVT U4898 ( .A1(n4999), .A2(n4854), .Y(n4986) );
  AND4X1_RVT U4899 ( .A1(n5000), .A2(n5001), .A3(n5002), .A4(n5003), .Y(n4999)
         );
  OR2X1_RVT U4900 ( .A1(n5004), .A2(n4819), .Y(n5002) );
  OR2X1_RVT U4901 ( .A1(n12692), .A2(n5005), .Y(n5001) );
  OR2X1_RVT U4902 ( .A1(n5006), .A2(n12700), .Y(n5000) );
  AND2X1_RVT U4903 ( .A1(n4897), .A2(n5007), .Y(n5006) );
  OR2X1_RVT U4904 ( .A1(n4899), .A2(n5008), .Y(n4985) );
  AND4X1_RVT U4905 ( .A1(n5009), .A2(n5010), .A3(n5011), .A4(n5012), .Y(n4917)
         );
  AND4X1_RVT U4906 ( .A1(n5013), .A2(n5014), .A3(n5015), .A4(n5016), .Y(n5012)
         );
  OR2X1_RVT U4907 ( .A1(n12696), .A2(n5017), .Y(n5016) );
  OR2X1_RVT U4908 ( .A1(n12697), .A2(n5018), .Y(n5015) );
  OR2X1_RVT U4909 ( .A1(n12694), .A2(n5019), .Y(n5014) );
  OR2X1_RVT U4910 ( .A1(n12444), .A2(n5020), .Y(n5013) );
  OR2X1_RVT U4911 ( .A1(n5021), .A2(n12451), .Y(n5010) );
  AND4X1_RVT U4912 ( .A1(n5023), .A2(n5024), .A3(n5025), .A4(n5026), .Y(n5022)
         );
  AND4X1_RVT U4913 ( .A1(n5027), .A2(n5028), .A3(n5029), .A4(n5030), .Y(n5026)
         );
  AND4X1_RVT U4914 ( .A1(n5031), .A2(n5032), .A3(n5033), .A4(n5034), .Y(n5030)
         );
  OR2X1_RVT U4915 ( .A1(n3168), .A2(n3969), .Y(n5034) );
  OR2X1_RVT U4916 ( .A1(n12883), .A2(n12503), .Y(n3969) );
  OR2X1_RVT U4917 ( .A1(n12477), .A2(n12487), .Y(n3168) );
  OR2X1_RVT U4918 ( .A1(n5035), .A2(n2754), .Y(n5033) );
  AND2X1_RVT U4919 ( .A1(n2700), .A2(n3924), .Y(n5035) );
  OR2X1_RVT U4920 ( .A1(n51), .A2(n5036), .Y(n2700) );
  OR2X1_RVT U4921 ( .A1(n12477), .A2(n12880), .Y(n5036) );
  OR2X1_RVT U4922 ( .A1(n5037), .A2(n2682), .Y(n5032) );
  OR2X1_RVT U4923 ( .A1(n12491), .A2(n2843), .Y(n2682) );
  AND2X1_RVT U4924 ( .A1(n2818), .A2(n5038), .Y(n5037) );
  OR2X1_RVT U4925 ( .A1(n2697), .A2(n2899), .Y(n5038) );
  OR2X1_RVT U4926 ( .A1(n12495), .A2(n12483), .Y(n2697) );
  OR2X1_RVT U4927 ( .A1(n2943), .A2(n5039), .Y(n2818) );
  OR2X1_RVT U4928 ( .A1(n12891), .A2(n12498), .Y(n5039) );
  OR2X1_RVT U4929 ( .A1(n5040), .A2(n2741), .Y(n5031) );
  AND2X1_RVT U4930 ( .A1(n3138), .A2(n5041), .Y(n5040) );
  OR2X1_RVT U4931 ( .A1(n5042), .A2(n12880), .Y(n5041) );
  AND2X1_RVT U4932 ( .A1(n2797), .A2(n3150), .Y(n5042) );
  OR2X1_RVT U4933 ( .A1(n12888), .A2(n2759), .Y(n3150) );
  OR2X1_RVT U4934 ( .A1(n12504), .A2(n5043), .Y(n3138) );
  OR2X1_RVT U4935 ( .A1(n12893), .A2(n12889), .Y(n5043) );
  OR2X1_RVT U4936 ( .A1(n5044), .A2(n12482), .Y(n5029) );
  AND2X1_RVT U4937 ( .A1(n5045), .A2(n5046), .Y(n5044) );
  OR2X1_RVT U4938 ( .A1(n5047), .A2(n2843), .Y(n5046) );
  AND2X1_RVT U4939 ( .A1(n2908), .A2(n5048), .Y(n5047) );
  OR2X1_RVT U4940 ( .A1(n2699), .A2(n2821), .Y(n5045) );
  OR2X1_RVT U4941 ( .A1(n12496), .A2(n2757), .Y(n2821) );
  OR2X1_RVT U4942 ( .A1(n5049), .A2(n12889), .Y(n5028) );
  AND2X1_RVT U4943 ( .A1(n2913), .A2(n3072), .Y(n5049) );
  OR2X1_RVT U4944 ( .A1(n12494), .A2(n5050), .Y(n3072) );
  OR2X1_RVT U4945 ( .A1(n2753), .A2(n12483), .Y(n5050) );
  OR2X1_RVT U4946 ( .A1(n2699), .A2(n3180), .Y(n2913) );
  OR2X1_RVT U4947 ( .A1(n12483), .A2(n12498), .Y(n3180) );
  OR2X1_RVT U4948 ( .A1(n5051), .A2(n12480), .Y(n5027) );
  AND2X1_RVT U4949 ( .A1(n2953), .A2(n5052), .Y(n5051) );
  OR2X1_RVT U4950 ( .A1(n3167), .A2(n2747), .Y(n5052) );
  OR2X1_RVT U4951 ( .A1(n2806), .A2(n3945), .Y(n2953) );
  OR2X1_RVT U4952 ( .A1(n12888), .A2(n51), .Y(n3945) );
  AND2X1_RVT U4953 ( .A1(n12484), .A2(n12891), .Y(n3049) );
  AND4X1_RVT U4954 ( .A1(n5053), .A2(n5054), .A3(n5055), .A4(n5056), .Y(n5025)
         );
  AND4X1_RVT U4955 ( .A1(n5057), .A2(n5058), .A3(n5059), .A4(n5060), .Y(n5056)
         );
  OR2X1_RVT U4956 ( .A1(n5061), .A2(n12489), .Y(n5060) );
  AND2X1_RVT U4957 ( .A1(n2940), .A2(n3011), .Y(n5061) );
  OR2X1_RVT U4958 ( .A1(n2756), .A2(n3924), .Y(n3011) );
  OR2X1_RVT U4959 ( .A1(n12891), .A2(n2753), .Y(n3924) );
  OR2X1_RVT U4960 ( .A1(n12878), .A2(n12479), .Y(n2756) );
  OR2X1_RVT U4961 ( .A1(n12480), .A2(n3043), .Y(n2940) );
  OR2X1_RVT U4962 ( .A1(n12484), .A2(n12498), .Y(n3043) );
  OR2X1_RVT U4963 ( .A1(n5062), .A2(n12887), .Y(n5059) );
  AND2X1_RVT U4964 ( .A1(n3102), .A2(n5063), .Y(n5062) );
  OR2X1_RVT U4965 ( .A1(n3060), .A2(n2770), .Y(n5063) );
  OR2X1_RVT U4966 ( .A1(n2943), .A2(n5064), .Y(n2770) );
  OR2X1_RVT U4967 ( .A1(n12509), .A2(n12485), .Y(n5064) );
  OR2X1_RVT U4968 ( .A1(n12493), .A2(n5065), .Y(n3102) );
  OR2X1_RVT U4969 ( .A1(n2943), .A2(n2739), .Y(n5065) );
  OR2X1_RVT U4970 ( .A1(n5066), .A2(n12893), .Y(n5058) );
  AND2X1_RVT U4971 ( .A1(n3048), .A2(n2977), .Y(n5066) );
  OR2X1_RVT U4972 ( .A1(n2759), .A2(n2795), .Y(n2977) );
  OR2X1_RVT U4973 ( .A1(n12885), .A2(n2943), .Y(n2795) );
  OR2X1_RVT U4974 ( .A1(n3167), .A2(n2775), .Y(n3048) );
  OR2X1_RVT U4975 ( .A1(n12490), .A2(n12890), .Y(n3167) );
  OR2X1_RVT U4976 ( .A1(n5067), .A2(n2817), .Y(n5057) );
  AND2X1_RVT U4977 ( .A1(n5068), .A2(n5069), .Y(n5067) );
  OR2X1_RVT U4978 ( .A1(n2739), .A2(n3166), .Y(n5069) );
  OR2X1_RVT U4979 ( .A1(n12887), .A2(n59), .Y(n3166) );
  AND2X1_RVT U4980 ( .A1(n5070), .A2(n3034), .Y(n5068) );
  OR2X1_RVT U4981 ( .A1(n2747), .A2(n5071), .Y(n3034) );
  OR2X1_RVT U4982 ( .A1(n12506), .A2(n12485), .Y(n5071) );
  OR2X1_RVT U4983 ( .A1(n2803), .A2(n2740), .Y(n5055) );
  OR2X1_RVT U4984 ( .A1(n12880), .A2(n2699), .Y(n2803) );
  OR2X1_RVT U4985 ( .A1(n5072), .A2(n2703), .Y(n5054) );
  AND2X1_RVT U4986 ( .A1(n5073), .A2(n2884), .Y(n5072) );
  AND2X1_RVT U4987 ( .A1(n5074), .A2(n5075), .Y(n2884) );
  OR2X1_RVT U4988 ( .A1(n12494), .A2(n2908), .Y(n5075) );
  OR2X1_RVT U4989 ( .A1(n2806), .A2(n2680), .Y(n5074) );
  OR2X1_RVT U4990 ( .A1(n12479), .A2(n2753), .Y(n2680) );
  AND2X1_RVT U4991 ( .A1(n5076), .A2(n3070), .Y(n5073) );
  OR2X1_RVT U4992 ( .A1(n2837), .A2(n3977), .Y(n3070) );
  OR2X1_RVT U4993 ( .A1(n12882), .A2(n49), .Y(n3977) );
  OR2X1_RVT U4994 ( .A1(n2699), .A2(n2866), .Y(n5076) );
  OR2X1_RVT U4995 ( .A1(n12478), .A2(n5077), .Y(n2866) );
  OR2X1_RVT U4996 ( .A1(n12878), .A2(n12507), .Y(n5077) );
  OR2X1_RVT U4997 ( .A1(n5078), .A2(n12878), .Y(n5053) );
  AND4X1_RVT U4998 ( .A1(n5079), .A2(n5080), .A3(n5081), .A4(n3212), .Y(n5078)
         );
  OR2X1_RVT U4999 ( .A1(n2753), .A2(n3133), .Y(n3212) );
  OR2X1_RVT U5000 ( .A1(n12883), .A2(n12889), .Y(n3133) );
  OR2X1_RVT U5001 ( .A1(n2753), .A2(n5082), .Y(n5081) );
  OR2X1_RVT U5002 ( .A1(n12484), .A2(n12489), .Y(n5082) );
  OR2X1_RVT U5003 ( .A1(n12888), .A2(n2712), .Y(n2753) );
  OR2X1_RVT U5004 ( .A1(n5083), .A2(n2834), .Y(n5080) );
  OR2X1_RVT U5005 ( .A1(n12478), .A2(n2678), .Y(n2834) );
  AND2X1_RVT U5006 ( .A1(n2817), .A2(n5084), .Y(n5083) );
  OR2X1_RVT U5007 ( .A1(n12886), .A2(n2717), .Y(n5084) );
  OR2X1_RVT U5008 ( .A1(n12882), .A2(n12489), .Y(n2817) );
  OR2X1_RVT U5009 ( .A1(n12884), .A2(n5048), .Y(n5079) );
  OR2X1_RVT U5010 ( .A1(n12888), .A2(n2757), .Y(n5048) );
  OR2X1_RVT U5011 ( .A1(n2703), .A2(n49), .Y(n2757) );
  AND4X1_RVT U5012 ( .A1(n5085), .A2(n5086), .A3(n5087), .A4(n5088), .Y(n5024)
         );
  AND4X1_RVT U5013 ( .A1(n5089), .A2(n5090), .A3(n5091), .A4(n5092), .Y(n5088)
         );
  OR2X1_RVT U5014 ( .A1(n2775), .A2(n2902), .Y(n5092) );
  OR2X1_RVT U5015 ( .A1(n12491), .A2(n2797), .Y(n2902) );
  OR2X1_RVT U5016 ( .A1(n12495), .A2(n2943), .Y(n2775) );
  OR2X1_RVT U5017 ( .A1(n2762), .A2(n3238), .Y(n5091) );
  OR2X1_RVT U5018 ( .A1(n12892), .A2(n12478), .Y(n3238) );
  OR2X1_RVT U5019 ( .A1(n2828), .A2(n2754), .Y(n2762) );
  OR2X1_RVT U5020 ( .A1(n2747), .A2(n2774), .Y(n5090) );
  OR2X1_RVT U5021 ( .A1(n12487), .A2(n12500), .Y(n2774) );
  OR2X1_RVT U5022 ( .A1(n12477), .A2(n12879), .Y(n2747) );
  OR2X1_RVT U5023 ( .A1(n59), .A2(n3113), .Y(n5089) );
  OR2X1_RVT U5024 ( .A1(n12485), .A2(n2900), .Y(n3113) );
  OR2X1_RVT U5025 ( .A1(n2717), .A2(n3147), .Y(n5087) );
  OR2X1_RVT U5026 ( .A1(n59), .A2(n5093), .Y(n3147) );
  OR2X1_RVT U5027 ( .A1(n12885), .A2(n12498), .Y(n5093) );
  AND2X1_RVT U5028 ( .A1(n12479), .A2(n12482), .Y(n3177) );
  OR2X1_RVT U5029 ( .A1(n2759), .A2(n2707), .Y(n5086) );
  OR2X1_RVT U5030 ( .A1(n12507), .A2(n5094), .Y(n2707) );
  OR2X1_RVT U5031 ( .A1(n12886), .A2(n12878), .Y(n5094) );
  OR2X1_RVT U5032 ( .A1(n12484), .A2(n2739), .Y(n2759) );
  OR2X1_RVT U5033 ( .A1(n2806), .A2(n5070), .Y(n5085) );
  OR2X1_RVT U5034 ( .A1(n12480), .A2(n2761), .Y(n5070) );
  OR2X1_RVT U5035 ( .A1(n12888), .A2(n12889), .Y(n2761) );
  AND4X1_RVT U5036 ( .A1(n5095), .A2(n2872), .A3(n5096), .A4(n5097), .Y(n5023)
         );
  OR2X1_RVT U5037 ( .A1(n12484), .A2(n3974), .Y(n5097) );
  OR2X1_RVT U5038 ( .A1(n12884), .A2(n2867), .Y(n3974) );
  OR2X1_RVT U5039 ( .A1(n12482), .A2(n2908), .Y(n2867) );
  OR2X1_RVT U5040 ( .A1(n12477), .A2(n2734), .Y(n2908) );
  AND2X1_RVT U5041 ( .A1(n5098), .A2(n5099), .Y(n5096) );
  OR2X1_RVT U5042 ( .A1(n12506), .A2(n3237), .Y(n5099) );
  OR2X1_RVT U5043 ( .A1(n2806), .A2(n2899), .Y(n3237) );
  OR2X1_RVT U5044 ( .A1(n12484), .A2(n12478), .Y(n2899) );
  OR2X1_RVT U5045 ( .A1(n12479), .A2(n2695), .Y(n2734) );
  OR2X1_RVT U5046 ( .A1(n12891), .A2(n2968), .Y(n5098) );
  OR2X1_RVT U5047 ( .A1(n12503), .A2(n3002), .Y(n2968) );
  OR2X1_RVT U5048 ( .A1(n12883), .A2(n12878), .Y(n3002) );
  OR2X1_RVT U5049 ( .A1(n12881), .A2(n12495), .Y(n2678) );
  AND2X1_RVT U5050 ( .A1(n5100), .A2(n5101), .Y(n2872) );
  OR2X1_RVT U5051 ( .A1(n2754), .A2(n2740), .Y(n5101) );
  OR2X1_RVT U5052 ( .A1(n12890), .A2(n2712), .Y(n2740) );
  AND2X1_RVT U5053 ( .A1(n2739), .A2(n2703), .Y(n2792) );
  OR2X1_RVT U5054 ( .A1(n12490), .A2(n2806), .Y(n2754) );
  OR2X1_RVT U5055 ( .A1(n12879), .A2(n2843), .Y(n2806) );
  OR2X1_RVT U5056 ( .A1(n5102), .A2(n2797), .Y(n5100) );
  OR2X1_RVT U5057 ( .A1(n12484), .A2(n49), .Y(n2797) );
  AND2X1_RVT U5058 ( .A1(n12892), .A2(n12477), .Y(n3060) );
  OR2X1_RVT U5059 ( .A1(n12483), .A2(n2900), .Y(n5102) );
  OR2X1_RVT U5060 ( .A1(n12888), .A2(n12500), .Y(n2900) );
  AND2X1_RVT U5061 ( .A1(n5103), .A2(n5104), .Y(n5095) );
  OR2X1_RVT U5062 ( .A1(n2720), .A2(n3053), .Y(n5104) );
  OR2X1_RVT U5063 ( .A1(n12485), .A2(n2760), .Y(n3053) );
  OR2X1_RVT U5064 ( .A1(n12500), .A2(n2837), .Y(n2760) );
  OR2X1_RVT U5065 ( .A1(n12480), .A2(n12483), .Y(n2837) );
  OR2X1_RVT U5066 ( .A1(n12885), .A2(n12883), .Y(n2699) );
  OR2X1_RVT U5067 ( .A1(n12893), .A2(n12887), .Y(n2720) );
  XOR2X1_RVT U5068 ( .A1(key[108]), .A2(state[108]), .Y(n2695) );
  OR2X1_RVT U5069 ( .A1(n2712), .A2(n2841), .Y(n5103) );
  OR2X1_RVT U5070 ( .A1(n2943), .A2(n3134), .Y(n2841) );
  OR2X1_RVT U5071 ( .A1(n12487), .A2(n2741), .Y(n3134) );
  OR2X1_RVT U5072 ( .A1(n12886), .A2(n2843), .Y(n2741) );
  XOR2X1_RVT U5073 ( .A1(key[106]), .A2(state[106]), .Y(n2843) );
  XOR2X1_RVT U5074 ( .A1(key[107]), .A2(state[107]), .Y(n2777) );
  OR2X1_RVT U5075 ( .A1(n12891), .A2(n12485), .Y(n2717) );
  XOR2X1_RVT U5076 ( .A1(key[109]), .A2(state[109]), .Y(n2703) );
  XOR2X1_RVT U5077 ( .A1(key[110]), .A2(state[110]), .Y(n2739) );
  OR2X1_RVT U5078 ( .A1(n12881), .A2(n12483), .Y(n2943) );
  XOR2X1_RVT U5079 ( .A1(key[104]), .A2(state[104]), .Y(n2718) );
  XOR2X1_RVT U5080 ( .A1(key[105]), .A2(state[105]), .Y(n2828) );
  XOR2X1_RVT U5081 ( .A1(key[111]), .A2(state[111]), .Y(n2712) );
  AND4X1_RVT U5082 ( .A1(n5106), .A2(n5107), .A3(n5108), .A4(n5109), .Y(n5105)
         );
  AND4X1_RVT U5083 ( .A1(n5110), .A2(n5111), .A3(n5112), .A4(n5113), .Y(n5109)
         );
  AND4X1_RVT U5084 ( .A1(n5114), .A2(n4808), .A3(n4978), .A4(n5115), .Y(n5113)
         );
  OR2X1_RVT U5085 ( .A1(n5116), .A2(n12691), .Y(n4808) );
  AND2X1_RVT U5086 ( .A1(n5117), .A2(n5118), .Y(n5116) );
  OR2X1_RVT U5087 ( .A1(n4852), .A2(n5119), .Y(n5118) );
  OR2X1_RVT U5088 ( .A1(n5120), .A2(n4934), .Y(n5117) );
  OR2X1_RVT U5089 ( .A1(n5121), .A2(n4893), .Y(n5114) );
  AND2X1_RVT U5090 ( .A1(n5122), .A2(n5123), .Y(n5121) );
  OR2X1_RVT U5091 ( .A1(n12696), .A2(n4877), .Y(n5123) );
  OR2X1_RVT U5092 ( .A1(n5124), .A2(n4836), .Y(n5112) );
  AND2X1_RVT U5093 ( .A1(n5125), .A2(n5126), .Y(n5124) );
  OR2X1_RVT U5094 ( .A1(n5127), .A2(n12702), .Y(n5126) );
  AND2X1_RVT U5095 ( .A1(n4884), .A2(n5128), .Y(n5127) );
  OR2X1_RVT U5096 ( .A1(n5129), .A2(n12471), .Y(n5111) );
  AND2X1_RVT U5097 ( .A1(n5130), .A2(n5131), .Y(n5129) );
  OR2X1_RVT U5098 ( .A1(n4877), .A2(n4843), .Y(n5131) );
  OR2X1_RVT U5099 ( .A1(n5132), .A2(n12454), .Y(n5110) );
  AND2X1_RVT U5100 ( .A1(n4961), .A2(n5133), .Y(n5132) );
  OR2X1_RVT U5101 ( .A1(n4890), .A2(n5134), .Y(n4961) );
  AND4X1_RVT U5102 ( .A1(n5135), .A2(n5136), .A3(n5137), .A4(n5138), .Y(n5108)
         );
  OR2X1_RVT U5103 ( .A1(n5139), .A2(n12461), .Y(n5138) );
  AND2X1_RVT U5104 ( .A1(n5140), .A2(n5141), .Y(n5139) );
  OR2X1_RVT U5105 ( .A1(n4934), .A2(n4834), .Y(n5141) );
  AND2X1_RVT U5106 ( .A1(n5142), .A2(n5143), .Y(n5140) );
  OR2X1_RVT U5107 ( .A1(n4974), .A2(n5119), .Y(n5142) );
  AND2X1_RVT U5108 ( .A1(n5144), .A2(n5145), .Y(n5137) );
  OR2X1_RVT U5109 ( .A1(n5146), .A2(n4965), .Y(n5145) );
  AND2X1_RVT U5110 ( .A1(n5147), .A2(n4873), .Y(n5146) );
  OR2X1_RVT U5111 ( .A1(n4819), .A2(n4934), .Y(n4873) );
  OR2X1_RVT U5112 ( .A1(n5148), .A2(n296), .Y(n5144) );
  AND2X1_RVT U5113 ( .A1(n5149), .A2(n5150), .Y(n5148) );
  OR2X1_RVT U5114 ( .A1(n5151), .A2(n12463), .Y(n5150) );
  AND2X1_RVT U5115 ( .A1(n5152), .A2(n5153), .Y(n5151) );
  OR2X1_RVT U5116 ( .A1(n12458), .A2(n4884), .Y(n5153) );
  OR2X1_RVT U5117 ( .A1(n12706), .A2(n12460), .Y(n5152) );
  AND2X1_RVT U5118 ( .A1(n4935), .A2(n5128), .Y(n5149) );
  OR2X1_RVT U5119 ( .A1(n4965), .A2(n5154), .Y(n4935) );
  OR2X1_RVT U5120 ( .A1(n12701), .A2(n12697), .Y(n5154) );
  OR2X1_RVT U5121 ( .A1(n5155), .A2(n4954), .Y(n5136) );
  AND4X1_RVT U5122 ( .A1(n4913), .A2(n5156), .A3(n5157), .A4(n5158), .Y(n5155)
         );
  OR2X1_RVT U5123 ( .A1(n12462), .A2(n4934), .Y(n5158) );
  AND2X1_RVT U5124 ( .A1(n5159), .A2(n5160), .Y(n5157) );
  OR2X1_RVT U5125 ( .A1(n12706), .A2(n12471), .Y(n5156) );
  AND2X1_RVT U5126 ( .A1(n5161), .A2(n5162), .Y(n4913) );
  OR2X1_RVT U5127 ( .A1(n5163), .A2(n294), .Y(n5162) );
  OR2X1_RVT U5128 ( .A1(n4877), .A2(n12691), .Y(n5161) );
  AND2X1_RVT U5129 ( .A1(n5164), .A2(n5165), .Y(n5135) );
  OR2X1_RVT U5130 ( .A1(n5166), .A2(n12693), .Y(n5165) );
  AND2X1_RVT U5131 ( .A1(n5167), .A2(n5168), .Y(n5166) );
  OR2X1_RVT U5132 ( .A1(n5169), .A2(n12465), .Y(n5168) );
  AND2X1_RVT U5133 ( .A1(n5170), .A2(n5171), .Y(n5169) );
  AND2X1_RVT U5134 ( .A1(n5172), .A2(n5173), .Y(n5167) );
  OR2X1_RVT U5135 ( .A1(n5174), .A2(n12474), .Y(n5164) );
  AND4X1_RVT U5136 ( .A1(n5175), .A2(n5176), .A3(n5177), .A4(n5178), .Y(n5174)
         );
  OR2X1_RVT U5137 ( .A1(n12705), .A2(n5179), .Y(n5177) );
  OR2X1_RVT U5138 ( .A1(n294), .A2(n4891), .Y(n5176) );
  OR2X1_RVT U5139 ( .A1(n4980), .A2(n4934), .Y(n5175) );
  AND4X1_RVT U5140 ( .A1(n5180), .A2(n5181), .A3(n5182), .A4(n5183), .Y(n5107)
         );
  AND2X1_RVT U5141 ( .A1(n5184), .A2(n4944), .Y(n5183) );
  OR2X1_RVT U5142 ( .A1(n12449), .A2(n4910), .Y(n4944) );
  AND2X1_RVT U5143 ( .A1(n5185), .A2(n5186), .Y(n5184) );
  OR2X1_RVT U5144 ( .A1(n5187), .A2(n4859), .Y(n5186) );
  OR2X1_RVT U5145 ( .A1(n4911), .A2(n4971), .Y(n5185) );
  OR2X1_RVT U5146 ( .A1(n294), .A2(n5188), .Y(n5182) );
  OR2X1_RVT U5147 ( .A1(n12704), .A2(n5189), .Y(n5181) );
  OR2X1_RVT U5148 ( .A1(n4980), .A2(n5190), .Y(n5180) );
  AND4X1_RVT U5149 ( .A1(n5191), .A2(n5192), .A3(n5193), .A4(n5194), .Y(n5106)
         );
  AND2X1_RVT U5150 ( .A1(n5195), .A2(n5196), .Y(n5194) );
  OR2X1_RVT U5151 ( .A1(n12444), .A2(n5197), .Y(n5196) );
  AND2X1_RVT U5152 ( .A1(n5198), .A2(n5199), .Y(n5195) );
  OR2X1_RVT U5153 ( .A1(n4876), .A2(n4886), .Y(n5199) );
  OR2X1_RVT U5154 ( .A1(n12465), .A2(n4936), .Y(n4886) );
  OR2X1_RVT U5155 ( .A1(n12451), .A2(n5200), .Y(n5198) );
  OR2X1_RVT U5156 ( .A1(n4857), .A2(n4850), .Y(n5193) );
  OR2X1_RVT U5157 ( .A1(n4943), .A2(n5201), .Y(n4850) );
  OR2X1_RVT U5158 ( .A1(n12700), .A2(n5202), .Y(n5192) );
  OR2X1_RVT U5159 ( .A1(n12463), .A2(n4977), .Y(n5191) );
  OR2X1_RVT U5160 ( .A1(n12691), .A2(n5122), .Y(n4977) );
  AND4X1_RVT U5161 ( .A1(n5204), .A2(n5205), .A3(n5206), .A4(n5207), .Y(n5203)
         );
  AND4X1_RVT U5162 ( .A1(n5208), .A2(n5209), .A3(n5210), .A4(n5211), .Y(n5207)
         );
  OR2X1_RVT U5163 ( .A1(n304), .A2(n5212), .Y(n5211) );
  OR2X1_RVT U5164 ( .A1(n5213), .A2(n12476), .Y(n5212) );
  AND2X1_RVT U5165 ( .A1(n12465), .A2(n4896), .Y(n5213) );
  AND2X1_RVT U5166 ( .A1(n4811), .A2(n5214), .Y(n5210) );
  OR2X1_RVT U5167 ( .A1(n12454), .A2(n5215), .Y(n4811) );
  OR2X1_RVT U5168 ( .A1(n304), .A2(n4890), .Y(n5215) );
  OR2X1_RVT U5169 ( .A1(n5216), .A2(n4819), .Y(n5209) );
  AND2X1_RVT U5170 ( .A1(n5217), .A2(n5218), .Y(n5216) );
  AND2X1_RVT U5171 ( .A1(n5219), .A2(n5220), .Y(n5208) );
  OR2X1_RVT U5172 ( .A1(n5221), .A2(n5222), .Y(n5220) );
  AND2X1_RVT U5173 ( .A1(n5223), .A2(n4900), .Y(n5221) );
  OR2X1_RVT U5174 ( .A1(n5224), .A2(n4891), .Y(n5219) );
  AND2X1_RVT U5175 ( .A1(n5159), .A2(n4910), .Y(n5224) );
  OR2X1_RVT U5176 ( .A1(n12452), .A2(n5225), .Y(n5159) );
  OR2X1_RVT U5177 ( .A1(n12706), .A2(n12462), .Y(n5225) );
  AND4X1_RVT U5178 ( .A1(n5226), .A2(n5227), .A3(n5228), .A4(n5229), .Y(n5206)
         );
  OR2X1_RVT U5179 ( .A1(n5230), .A2(n12696), .Y(n5229) );
  AND2X1_RVT U5180 ( .A1(n4959), .A2(n5231), .Y(n5230) );
  OR2X1_RVT U5181 ( .A1(n12704), .A2(n5004), .Y(n4959) );
  AND2X1_RVT U5182 ( .A1(n5232), .A2(n5233), .Y(n5228) );
  OR2X1_RVT U5183 ( .A1(n5234), .A2(n12694), .Y(n5233) );
  AND2X1_RVT U5184 ( .A1(n5235), .A2(n5236), .Y(n5234) );
  OR2X1_RVT U5185 ( .A1(n4854), .A2(n5179), .Y(n5236) );
  OR2X1_RVT U5186 ( .A1(n5237), .A2(n12692), .Y(n5232) );
  AND2X1_RVT U5187 ( .A1(n5238), .A2(n5239), .Y(n5237) );
  OR2X1_RVT U5188 ( .A1(n5240), .A2(n12465), .Y(n5227) );
  AND2X1_RVT U5189 ( .A1(n5241), .A2(n5242), .Y(n5240) );
  AND2X1_RVT U5190 ( .A1(n5243), .A2(n5244), .Y(n5241) );
  AND2X1_RVT U5191 ( .A1(n5245), .A2(n5246), .Y(n5226) );
  OR2X1_RVT U5192 ( .A1(n5247), .A2(n5163), .Y(n5246) );
  AND2X1_RVT U5193 ( .A1(n5248), .A2(n4911), .Y(n5247) );
  AND2X1_RVT U5194 ( .A1(n5249), .A2(n5250), .Y(n5248) );
  OR2X1_RVT U5195 ( .A1(n5251), .A2(n12468), .Y(n5245) );
  AND2X1_RVT U5196 ( .A1(n5252), .A2(n5253), .Y(n5251) );
  OR2X1_RVT U5197 ( .A1(n12703), .A2(n12470), .Y(n5253) );
  AND2X1_RVT U5198 ( .A1(n4900), .A2(n5254), .Y(n5252) );
  AND4X1_RVT U5199 ( .A1(n5255), .A2(n5256), .A3(n5257), .A4(n5258), .Y(n5205)
         );
  AND2X1_RVT U5200 ( .A1(n5259), .A2(n5260), .Y(n5258) );
  OR2X1_RVT U5201 ( .A1(n4893), .A2(n4967), .Y(n5260) );
  OR2X1_RVT U5202 ( .A1(n12698), .A2(n4900), .Y(n4967) );
  AND2X1_RVT U5203 ( .A1(n5261), .A2(n5262), .Y(n5259) );
  OR2X1_RVT U5204 ( .A1(n5128), .A2(n4859), .Y(n5262) );
  OR2X1_RVT U5205 ( .A1(n12705), .A2(n12461), .Y(n4859) );
  OR2X1_RVT U5206 ( .A1(n4943), .A2(n4993), .Y(n5261) );
  OR2X1_RVT U5207 ( .A1(n12693), .A2(n5263), .Y(n4993) );
  OR2X1_RVT U5208 ( .A1(n5264), .A2(n12444), .Y(n5257) );
  AND4X1_RVT U5209 ( .A1(n5265), .A2(n5266), .A3(n5267), .A4(n5268), .Y(n5264)
         );
  OR2X1_RVT U5210 ( .A1(n5201), .A2(n4891), .Y(n5267) );
  OR2X1_RVT U5211 ( .A1(n5269), .A2(n4888), .Y(n5266) );
  OR2X1_RVT U5212 ( .A1(n12702), .A2(n4843), .Y(n5265) );
  OR2X1_RVT U5213 ( .A1(n5270), .A2(n12445), .Y(n5256) );
  AND2X1_RVT U5214 ( .A1(n5271), .A2(n5272), .Y(n5270) );
  OR2X1_RVT U5215 ( .A1(n5201), .A2(n4843), .Y(n5272) );
  AND2X1_RVT U5216 ( .A1(n5273), .A2(n5202), .Y(n5271) );
  OR2X1_RVT U5217 ( .A1(n4891), .A2(n5274), .Y(n5202) );
  OR2X1_RVT U5218 ( .A1(n12693), .A2(n12705), .Y(n5274) );
  OR2X1_RVT U5219 ( .A1(n5275), .A2(n12452), .Y(n5255) );
  AND4X1_RVT U5220 ( .A1(n5276), .A2(n5189), .A3(n4915), .A4(n4887), .Y(n5275)
         );
  OR2X1_RVT U5221 ( .A1(n4912), .A2(n5277), .Y(n4887) );
  OR2X1_RVT U5222 ( .A1(n12695), .A2(n4849), .Y(n5277) );
  OR2X1_RVT U5223 ( .A1(n4974), .A2(n5008), .Y(n4915) );
  OR2X1_RVT U5224 ( .A1(n4893), .A2(n5278), .Y(n5189) );
  OR2X1_RVT U5225 ( .A1(n12476), .A2(n12445), .Y(n5278) );
  OR2X1_RVT U5226 ( .A1(n4852), .A2(n5279), .Y(n5276) );
  OR2X1_RVT U5227 ( .A1(n5280), .A2(n12450), .Y(n5279) );
  AND4X1_RVT U5228 ( .A1(n5281), .A2(n5282), .A3(n5283), .A4(n5284), .Y(n5204)
         );
  AND2X1_RVT U5229 ( .A1(n5285), .A2(n5286), .Y(n5284) );
  AND2X1_RVT U5230 ( .A1(n5287), .A2(n5288), .Y(n5285) );
  OR2X1_RVT U5231 ( .A1(n4884), .A2(n5242), .Y(n5288) );
  OR2X1_RVT U5232 ( .A1(n4896), .A2(n5289), .Y(n5242) );
  OR2X1_RVT U5233 ( .A1(n12694), .A2(n12696), .Y(n5289) );
  OR2X1_RVT U5234 ( .A1(n12701), .A2(n5290), .Y(n5287) );
  OR2X1_RVT U5235 ( .A1(n12461), .A2(n5291), .Y(n5283) );
  OR2X1_RVT U5236 ( .A1(n12704), .A2(n5292), .Y(n5282) );
  OR2X1_RVT U5237 ( .A1(n4896), .A2(n5293), .Y(n5281) );
  AND4X1_RVT U5238 ( .A1(n5295), .A2(n5296), .A3(n5297), .A4(n5298), .Y(n5294)
         );
  AND4X1_RVT U5239 ( .A1(n5299), .A2(n5300), .A3(n5301), .A4(n5302), .Y(n5298)
         );
  AND4X1_RVT U5240 ( .A1(n5303), .A2(n5304), .A3(n4813), .A4(n5305), .Y(n5302)
         );
  OR2X1_RVT U5241 ( .A1(n4954), .A2(n5306), .Y(n4813) );
  OR2X1_RVT U5242 ( .A1(n5128), .A2(n296), .Y(n5306) );
  OR2X1_RVT U5243 ( .A1(n4817), .A2(n5307), .Y(n5304) );
  OR2X1_RVT U5244 ( .A1(n12699), .A2(n12702), .Y(n5307) );
  OR2X1_RVT U5245 ( .A1(n5163), .A2(n5308), .Y(n5303) );
  OR2X1_RVT U5246 ( .A1(n5309), .A2(n4854), .Y(n5308) );
  AND2X1_RVT U5247 ( .A1(n12465), .A2(n4954), .Y(n5309) );
  OR2X1_RVT U5248 ( .A1(n5310), .A2(n12471), .Y(n5301) );
  AND2X1_RVT U5249 ( .A1(n5178), .A2(n5250), .Y(n5310) );
  OR2X1_RVT U5250 ( .A1(n296), .A2(n5311), .Y(n5250) );
  OR2X1_RVT U5251 ( .A1(n12444), .A2(n12698), .Y(n5311) );
  OR2X1_RVT U5252 ( .A1(n4884), .A2(n5312), .Y(n5178) );
  OR2X1_RVT U5253 ( .A1(n12696), .A2(n4876), .Y(n5312) );
  OR2X1_RVT U5254 ( .A1(n5313), .A2(n4834), .Y(n5300) );
  AND2X1_RVT U5255 ( .A1(n5314), .A2(n5122), .Y(n5313) );
  OR2X1_RVT U5256 ( .A1(n4940), .A2(n4934), .Y(n5299) );
  AND4X1_RVT U5257 ( .A1(n5315), .A2(n5316), .A3(n5317), .A4(n5318), .Y(n5297)
         );
  AND2X1_RVT U5258 ( .A1(n5319), .A2(n5320), .Y(n5318) );
  OR2X1_RVT U5259 ( .A1(n5321), .A2(n12465), .Y(n5320) );
  AND2X1_RVT U5260 ( .A1(n5322), .A2(n4907), .Y(n5321) );
  AND2X1_RVT U5261 ( .A1(n5323), .A2(n5324), .Y(n5319) );
  OR2X1_RVT U5262 ( .A1(n5325), .A2(n4890), .Y(n5324) );
  AND2X1_RVT U5263 ( .A1(n4861), .A2(n4833), .Y(n5325) );
  OR2X1_RVT U5264 ( .A1(n12704), .A2(n4932), .Y(n4861) );
  OR2X1_RVT U5265 ( .A1(n5326), .A2(n4943), .Y(n5323) );
  AND2X1_RVT U5266 ( .A1(n5218), .A2(n5327), .Y(n5326) );
  OR2X1_RVT U5267 ( .A1(n12705), .A2(n4971), .Y(n5218) );
  OR2X1_RVT U5268 ( .A1(n5328), .A2(n12696), .Y(n5317) );
  AND2X1_RVT U5269 ( .A1(n4838), .A2(n5329), .Y(n5328) );
  OR2X1_RVT U5270 ( .A1(n4974), .A2(n4898), .Y(n5329) );
  OR2X1_RVT U5271 ( .A1(n4877), .A2(n5163), .Y(n4838) );
  OR2X1_RVT U5272 ( .A1(n5330), .A2(n294), .Y(n5316) );
  AND2X1_RVT U5273 ( .A1(n4888), .A2(n5331), .Y(n5330) );
  OR2X1_RVT U5274 ( .A1(n5332), .A2(n12449), .Y(n5331) );
  AND2X1_RVT U5275 ( .A1(n5333), .A2(n5334), .Y(n5332) );
  OR2X1_RVT U5276 ( .A1(n12697), .A2(n4871), .Y(n5334) );
  OR2X1_RVT U5277 ( .A1(n12476), .A2(n4974), .Y(n4888) );
  OR2X1_RVT U5278 ( .A1(n5335), .A2(n4958), .Y(n5315) );
  AND2X1_RVT U5279 ( .A1(n4891), .A2(n4936), .Y(n5335) );
  OR2X1_RVT U5280 ( .A1(n12693), .A2(n4819), .Y(n4936) );
  AND4X1_RVT U5281 ( .A1(n5336), .A2(n5337), .A3(n5338), .A4(n5339), .Y(n5296)
         );
  AND4X1_RVT U5282 ( .A1(n5340), .A2(n5341), .A3(n5342), .A4(n5343), .Y(n5339)
         );
  OR2X1_RVT U5283 ( .A1(n5344), .A2(n12704), .Y(n5343) );
  AND2X1_RVT U5284 ( .A1(n4994), .A2(n5345), .Y(n5344) );
  OR2X1_RVT U5285 ( .A1(n12473), .A2(n4843), .Y(n5345) );
  OR2X1_RVT U5286 ( .A1(n5346), .A2(n4836), .Y(n5342) );
  AND2X1_RVT U5287 ( .A1(n5347), .A2(n5348), .Y(n5346) );
  OR2X1_RVT U5288 ( .A1(n5349), .A2(n4871), .Y(n5348) );
  AND2X1_RVT U5289 ( .A1(n4896), .A2(n4884), .Y(n5349) );
  AND2X1_RVT U5290 ( .A1(n4898), .A2(n5223), .Y(n5347) );
  OR2X1_RVT U5291 ( .A1(n12474), .A2(n5119), .Y(n5223) );
  OR2X1_RVT U5292 ( .A1(n5350), .A2(n12463), .Y(n5341) );
  AND2X1_RVT U5293 ( .A1(n5351), .A2(n5352), .Y(n5350) );
  OR2X1_RVT U5294 ( .A1(n4884), .A2(n5353), .Y(n5352) );
  AND2X1_RVT U5295 ( .A1(n4966), .A2(n5243), .Y(n5351) );
  OR2X1_RVT U5296 ( .A1(n4876), .A2(n5134), .Y(n5243) );
  OR2X1_RVT U5297 ( .A1(n4849), .A2(n5354), .Y(n4966) );
  OR2X1_RVT U5298 ( .A1(n5355), .A2(n4819), .Y(n5340) );
  AND4X1_RVT U5299 ( .A1(n5356), .A2(n5357), .A3(n5358), .A4(n5291), .Y(n5355)
         );
  OR2X1_RVT U5300 ( .A1(n4912), .A2(n5359), .Y(n5291) );
  OR2X1_RVT U5301 ( .A1(n12444), .A2(n4876), .Y(n5359) );
  OR2X1_RVT U5302 ( .A1(n12701), .A2(n5201), .Y(n5357) );
  OR2X1_RVT U5303 ( .A1(n4877), .A2(n4974), .Y(n5356) );
  OR2X1_RVT U5304 ( .A1(n5128), .A2(n5170), .Y(n5338) );
  OR2X1_RVT U5305 ( .A1(n5360), .A2(n12447), .Y(n5337) );
  AND4X1_RVT U5306 ( .A1(n5361), .A2(n5362), .A3(n4921), .A4(n5019), .Y(n5360)
         );
  OR2X1_RVT U5307 ( .A1(n4843), .A2(n5008), .Y(n5019) );
  OR2X1_RVT U5308 ( .A1(n12701), .A2(n294), .Y(n5008) );
  OR2X1_RVT U5309 ( .A1(n4836), .A2(n4900), .Y(n4921) );
  OR2X1_RVT U5310 ( .A1(n12693), .A2(n5354), .Y(n5336) );
  AND4X1_RVT U5311 ( .A1(n5363), .A2(n5364), .A3(n5365), .A4(n5366), .Y(n5295)
         );
  OR2X1_RVT U5312 ( .A1(n12452), .A2(n5367), .Y(n5366) );
  AND2X1_RVT U5313 ( .A1(n5368), .A2(n5369), .Y(n5365) );
  OR2X1_RVT U5314 ( .A1(n12473), .A2(n5122), .Y(n5369) );
  OR2X1_RVT U5315 ( .A1(n4826), .A2(n4900), .Y(n5368) );
  OR2X1_RVT U5316 ( .A1(n296), .A2(n4857), .Y(n4900) );
  OR2X1_RVT U5317 ( .A1(n12476), .A2(n5018), .Y(n5364) );
  OR2X1_RVT U5318 ( .A1(n4893), .A2(n5370), .Y(n5018) );
  AND2X1_RVT U5319 ( .A1(n5371), .A2(n5372), .Y(n5363) );
  OR2X1_RVT U5320 ( .A1(n12445), .A2(n5373), .Y(n5372) );
  OR2X1_RVT U5321 ( .A1(n4896), .A2(n4845), .Y(n5371) );
  OR2X1_RVT U5322 ( .A1(n4819), .A2(n5187), .Y(n4845) );
  AND4X1_RVT U5323 ( .A1(n5375), .A2(n5376), .A3(n5377), .A4(n5378), .Y(n5374)
         );
  AND4X1_RVT U5324 ( .A1(n5379), .A2(n5380), .A3(n5381), .A4(n5382), .Y(n5378)
         );
  AND4X1_RVT U5325 ( .A1(n5115), .A2(n5305), .A3(n5383), .A4(n5384), .Y(n5382)
         );
  OR2X1_RVT U5326 ( .A1(n5385), .A2(n5386), .Y(n5305) );
  OR2X1_RVT U5327 ( .A1(n4817), .A2(n5170), .Y(n5115) );
  OR2X1_RVT U5328 ( .A1(n12702), .A2(n12461), .Y(n5170) );
  AND4X1_RVT U5329 ( .A1(n5373), .A2(n5239), .A3(n5362), .A4(n4814), .Y(n5381)
         );
  OR2X1_RVT U5330 ( .A1(n5387), .A2(n5004), .Y(n4814) );
  OR2X1_RVT U5331 ( .A1(n4819), .A2(n5388), .Y(n5362) );
  OR2X1_RVT U5332 ( .A1(n4852), .A2(n294), .Y(n5239) );
  OR2X1_RVT U5333 ( .A1(n4843), .A2(n5389), .Y(n5373) );
  OR2X1_RVT U5334 ( .A1(n12451), .A2(n12471), .Y(n5389) );
  AND4X1_RVT U5335 ( .A1(n5390), .A2(n5391), .A3(n5392), .A4(n5393), .Y(n5380)
         );
  OR2X1_RVT U5336 ( .A1(n5179), .A2(n5394), .Y(n5393) );
  OR2X1_RVT U5337 ( .A1(n12471), .A2(n4876), .Y(n5394) );
  OR2X1_RVT U5338 ( .A1(n5005), .A2(n5395), .Y(n5392) );
  OR2X1_RVT U5339 ( .A1(n12703), .A2(n4893), .Y(n5395) );
  OR2X1_RVT U5340 ( .A1(n5314), .A2(n5396), .Y(n5391) );
  OR2X1_RVT U5341 ( .A1(n5397), .A2(n4890), .Y(n5396) );
  OR2X1_RVT U5342 ( .A1(n12468), .A2(n5398), .Y(n5390) );
  OR2X1_RVT U5343 ( .A1(n5399), .A2(n12451), .Y(n5398) );
  AND2X1_RVT U5344 ( .A1(n5187), .A2(n5400), .Y(n5399) );
  AND2X1_RVT U5345 ( .A1(n5401), .A2(n5402), .Y(n5379) );
  OR2X1_RVT U5346 ( .A1(n5403), .A2(n4871), .Y(n5402) );
  AND2X1_RVT U5347 ( .A1(n5404), .A2(n5405), .Y(n5403) );
  OR2X1_RVT U5348 ( .A1(n12450), .A2(n5147), .Y(n5405) );
  OR2X1_RVT U5349 ( .A1(n12454), .A2(n5222), .Y(n5404) );
  AND2X1_RVT U5350 ( .A1(n5406), .A2(n5407), .Y(n5401) );
  OR2X1_RVT U5351 ( .A1(n5408), .A2(n4910), .Y(n5407) );
  AND2X1_RVT U5352 ( .A1(n5409), .A2(n5410), .Y(n5408) );
  OR2X1_RVT U5353 ( .A1(n12457), .A2(n304), .Y(n5410) );
  NAND2X1_RVT U5354 ( .A1(n4893), .A2(n12695), .Y(n5409) );
  OR2X1_RVT U5355 ( .A1(n5411), .A2(n296), .Y(n5406) );
  AND2X1_RVT U5356 ( .A1(n5200), .A2(n4994), .Y(n5411) );
  OR2X1_RVT U5357 ( .A1(n4843), .A2(n5412), .Y(n4994) );
  OR2X1_RVT U5358 ( .A1(n12706), .A2(n12446), .Y(n5412) );
  AND4X1_RVT U5359 ( .A1(n5011), .A2(n5413), .A3(n5286), .A4(n5414), .Y(n5377)
         );
  AND4X1_RVT U5360 ( .A1(n5415), .A2(n5416), .A3(n5417), .A4(n5418), .Y(n5414)
         );
  OR2X1_RVT U5361 ( .A1(n4974), .A2(n4895), .Y(n5418) );
  OR2X1_RVT U5362 ( .A1(n4912), .A2(n4941), .Y(n5417) );
  OR2X1_RVT U5363 ( .A1(n12694), .A2(n5249), .Y(n5416) );
  OR2X1_RVT U5364 ( .A1(n4890), .A2(n4872), .Y(n5249) );
  OR2X1_RVT U5365 ( .A1(n12702), .A2(n4954), .Y(n4872) );
  OR2X1_RVT U5366 ( .A1(n12460), .A2(n4995), .Y(n5415) );
  OR2X1_RVT U5367 ( .A1(n4876), .A2(n5187), .Y(n4995) );
  OR2X1_RVT U5368 ( .A1(n12444), .A2(n5163), .Y(n5187) );
  AND2X1_RVT U5369 ( .A1(n5419), .A2(n5420), .Y(n5286) );
  OR2X1_RVT U5370 ( .A1(n5421), .A2(n4943), .Y(n5420) );
  OR2X1_RVT U5371 ( .A1(n12470), .A2(n296), .Y(n5421) );
  OR2X1_RVT U5372 ( .A1(n5422), .A2(n4826), .Y(n5419) );
  OR2X1_RVT U5373 ( .A1(n12693), .A2(n4943), .Y(n4826) );
  OR2X1_RVT U5374 ( .A1(n4840), .A2(n4890), .Y(n5422) );
  OR2X1_RVT U5375 ( .A1(n12452), .A2(n5292), .Y(n5413) );
  AND2X1_RVT U5376 ( .A1(n5423), .A2(n5424), .Y(n5011) );
  OR2X1_RVT U5377 ( .A1(n4894), .A2(n4932), .Y(n5424) );
  OR2X1_RVT U5378 ( .A1(n5425), .A2(n5426), .Y(n5423) );
  AND4X1_RVT U5379 ( .A1(n5427), .A2(n5428), .A3(n5429), .A4(n5430), .Y(n5376)
         );
  OR2X1_RVT U5380 ( .A1(n5431), .A2(n5163), .Y(n5430) );
  AND2X1_RVT U5381 ( .A1(n5432), .A2(n5172), .Y(n5431) );
  OR2X1_RVT U5382 ( .A1(n12458), .A2(n5388), .Y(n5172) );
  OR2X1_RVT U5383 ( .A1(n5433), .A2(n12699), .Y(n5429) );
  AND2X1_RVT U5384 ( .A1(n5017), .A2(n4982), .Y(n5433) );
  OR2X1_RVT U5385 ( .A1(n12693), .A2(n4958), .Y(n4982) );
  OR2X1_RVT U5386 ( .A1(n5434), .A2(n5120), .Y(n5428) );
  AND2X1_RVT U5387 ( .A1(n5435), .A2(n5436), .Y(n5434) );
  OR2X1_RVT U5388 ( .A1(n12447), .A2(n4896), .Y(n5436) );
  AND2X1_RVT U5389 ( .A1(n5437), .A2(n4934), .Y(n5435) );
  OR2X1_RVT U5390 ( .A1(n294), .A2(n4893), .Y(n5437) );
  OR2X1_RVT U5391 ( .A1(n5438), .A2(n4834), .Y(n5427) );
  AND2X1_RVT U5392 ( .A1(n5439), .A2(n5440), .Y(n5438) );
  NAND2X1_RVT U5393 ( .A1(n4819), .A2(n5280), .Y(n5440) );
  AND2X1_RVT U5394 ( .A1(n5441), .A2(n5130), .Y(n5439) );
  OR2X1_RVT U5395 ( .A1(n4980), .A2(n5388), .Y(n5130) );
  OR2X1_RVT U5396 ( .A1(n12467), .A2(n5442), .Y(n5441) );
  AND4X1_RVT U5397 ( .A1(n5443), .A2(n5444), .A3(n5445), .A4(n5446), .Y(n5375)
         );
  OR2X1_RVT U5398 ( .A1(n5447), .A2(n4857), .Y(n5446) );
  AND2X1_RVT U5399 ( .A1(n5448), .A2(n4998), .Y(n5447) );
  AND2X1_RVT U5400 ( .A1(n5449), .A2(n5020), .Y(n5448) );
  OR2X1_RVT U5401 ( .A1(n296), .A2(n5426), .Y(n5020) );
  OR2X1_RVT U5402 ( .A1(n12446), .A2(n4954), .Y(n5426) );
  OR2X1_RVT U5403 ( .A1(n5450), .A2(n12463), .Y(n5445) );
  AND2X1_RVT U5404 ( .A1(n5451), .A2(n5452), .Y(n5450) );
  OR2X1_RVT U5405 ( .A1(n5453), .A2(n12691), .Y(n5452) );
  AND2X1_RVT U5406 ( .A1(n5454), .A2(n5455), .Y(n5453) );
  OR2X1_RVT U5407 ( .A1(n12445), .A2(n5314), .Y(n5455) );
  OR2X1_RVT U5408 ( .A1(n12698), .A2(n4877), .Y(n5454) );
  AND2X1_RVT U5409 ( .A1(n5456), .A2(n5457), .Y(n5451) );
  OR2X1_RVT U5410 ( .A1(n4843), .A2(n5458), .Y(n5456) );
  OR2X1_RVT U5411 ( .A1(n5459), .A2(n4877), .Y(n5444) );
  AND4X1_RVT U5412 ( .A1(n5460), .A2(n5461), .A3(n5462), .A4(n4843), .Y(n5459)
         );
  OR2X1_RVT U5413 ( .A1(n12699), .A2(n4893), .Y(n5462) );
  OR2X1_RVT U5414 ( .A1(n12457), .A2(n4912), .Y(n5461) );
  OR2X1_RVT U5415 ( .A1(n4965), .A2(n4943), .Y(n5460) );
  OR2X1_RVT U5416 ( .A1(n5463), .A2(n4819), .Y(n5443) );
  AND4X1_RVT U5417 ( .A1(n5327), .A2(n5464), .A3(n5125), .A4(n4958), .Y(n5463)
         );
  OR2X1_RVT U5418 ( .A1(n4912), .A2(n5458), .Y(n5125) );
  OR2X1_RVT U5419 ( .A1(n5163), .A2(n5370), .Y(n5464) );
  OR2X1_RVT U5420 ( .A1(n12451), .A2(n5128), .Y(n5327) );
  AND4X1_RVT U5421 ( .A1(n5466), .A2(n5467), .A3(n5468), .A4(n5469), .Y(n5465)
         );
  AND4X1_RVT U5422 ( .A1(n4895), .A2(n5214), .A3(n5470), .A4(n5471), .Y(n5469)
         );
  AND4X1_RVT U5423 ( .A1(n5293), .A2(n5238), .A3(n5383), .A4(n5384), .Y(n5471)
         );
  OR2X1_RVT U5424 ( .A1(n5386), .A2(n4816), .Y(n5384) );
  OR2X1_RVT U5425 ( .A1(n12697), .A2(n4934), .Y(n4816) );
  OR2X1_RVT U5426 ( .A1(n4833), .A2(n5425), .Y(n5383) );
  OR2X1_RVT U5427 ( .A1(n12702), .A2(n12465), .Y(n5425) );
  OR2X1_RVT U5428 ( .A1(n12691), .A2(n4954), .Y(n4833) );
  OR2X1_RVT U5429 ( .A1(n12703), .A2(n4852), .Y(n5238) );
  OR2X1_RVT U5430 ( .A1(n12474), .A2(n12458), .Y(n4852) );
  OR2X1_RVT U5431 ( .A1(n4974), .A2(n5472), .Y(n5293) );
  OR2X1_RVT U5432 ( .A1(n12465), .A2(n4878), .Y(n5472) );
  OR2X1_RVT U5433 ( .A1(n4876), .A2(n5473), .Y(n5470) );
  OR2X1_RVT U5434 ( .A1(n5004), .A2(n12456), .Y(n5473) );
  OR2X1_RVT U5435 ( .A1(n4943), .A2(n5474), .Y(n5214) );
  OR2X1_RVT U5436 ( .A1(n4877), .A2(n12463), .Y(n5474) );
  OR2X1_RVT U5437 ( .A1(n12695), .A2(n5385), .Y(n4895) );
  OR2X1_RVT U5438 ( .A1(n12458), .A2(n4894), .Y(n5385) );
  AND4X1_RVT U5439 ( .A1(n5475), .A2(n5476), .A3(n5477), .A4(n5478), .Y(n5468)
         );
  AND4X1_RVT U5440 ( .A1(n5479), .A2(n5480), .A3(n5481), .A4(n5482), .Y(n5478)
         );
  OR2X1_RVT U5441 ( .A1(n4910), .A2(n5483), .Y(n5482) );
  OR2X1_RVT U5442 ( .A1(n12447), .A2(n4980), .Y(n5483) );
  OR2X1_RVT U5443 ( .A1(n4893), .A2(n5484), .Y(n5481) );
  OR2X1_RVT U5444 ( .A1(n5485), .A2(n4857), .Y(n5484) );
  AND2X1_RVT U5445 ( .A1(n4836), .A2(n4896), .Y(n5485) );
  OR2X1_RVT U5446 ( .A1(n5486), .A2(n5487), .Y(n5480) );
  AND2X1_RVT U5447 ( .A1(n5134), .A2(n5007), .Y(n5486) );
  OR2X1_RVT U5448 ( .A1(n12696), .A2(n304), .Y(n5007) );
  OR2X1_RVT U5449 ( .A1(n12692), .A2(n12468), .Y(n5134) );
  OR2X1_RVT U5450 ( .A1(n5488), .A2(n4891), .Y(n5479) );
  AND2X1_RVT U5451 ( .A1(n5370), .A2(n5489), .Y(n5488) );
  OR2X1_RVT U5452 ( .A1(n12694), .A2(n296), .Y(n5489) );
  OR2X1_RVT U5453 ( .A1(n5490), .A2(n12470), .Y(n5477) );
  AND2X1_RVT U5454 ( .A1(n5361), .A2(n5491), .Y(n5490) );
  OR2X1_RVT U5455 ( .A1(n4884), .A2(n5314), .Y(n5491) );
  OR2X1_RVT U5456 ( .A1(n12451), .A2(n5179), .Y(n5361) );
  OR2X1_RVT U5457 ( .A1(n12698), .A2(n4884), .Y(n5179) );
  OR2X1_RVT U5458 ( .A1(n5492), .A2(n5128), .Y(n5476) );
  AND2X1_RVT U5459 ( .A1(n4998), .A2(n5353), .Y(n5492) );
  OR2X1_RVT U5460 ( .A1(n4854), .A2(n4943), .Y(n4998) );
  OR2X1_RVT U5461 ( .A1(n5493), .A2(n4934), .Y(n5475) );
  AND2X1_RVT U5462 ( .A1(n4897), .A2(n4899), .Y(n5493) );
  AND4X1_RVT U5463 ( .A1(n5494), .A2(n5495), .A3(n5496), .A4(n5497), .Y(n5467)
         );
  AND4X1_RVT U5464 ( .A1(n5498), .A2(n5499), .A3(n5500), .A4(n5501), .Y(n5497)
         );
  OR2X1_RVT U5465 ( .A1(n5502), .A2(n12454), .Y(n5501) );
  AND2X1_RVT U5466 ( .A1(n4825), .A2(n5200), .Y(n5502) );
  OR2X1_RVT U5467 ( .A1(n4974), .A2(n5005), .Y(n5200) );
  OR2X1_RVT U5468 ( .A1(n12457), .A2(n4857), .Y(n5005) );
  OR2X1_RVT U5469 ( .A1(n12461), .A2(n5503), .Y(n4825) );
  OR2X1_RVT U5470 ( .A1(n12444), .A2(n12450), .Y(n5503) );
  OR2X1_RVT U5471 ( .A1(n5504), .A2(n12468), .Y(n5500) );
  AND2X1_RVT U5472 ( .A1(n5217), .A2(n5505), .Y(n5504) );
  OR2X1_RVT U5473 ( .A1(n12473), .A2(n294), .Y(n5505) );
  OR2X1_RVT U5474 ( .A1(n12471), .A2(n4941), .Y(n5217) );
  OR2X1_RVT U5475 ( .A1(n5506), .A2(n12449), .Y(n5499) );
  AND2X1_RVT U5476 ( .A1(n5235), .A2(n5507), .Y(n5506) );
  OR2X1_RVT U5477 ( .A1(n12474), .A2(n4877), .Y(n5507) );
  OR2X1_RVT U5478 ( .A1(n4819), .A2(n5508), .Y(n5235) );
  OR2X1_RVT U5479 ( .A1(n5509), .A2(n4878), .Y(n5498) );
  AND2X1_RVT U5480 ( .A1(n5510), .A2(n5511), .Y(n5509) );
  OR2X1_RVT U5481 ( .A1(n4934), .A2(n12471), .Y(n5511) );
  AND2X1_RVT U5482 ( .A1(n5512), .A2(n4910), .Y(n5510) );
  OR2X1_RVT U5483 ( .A1(n4896), .A2(n4857), .Y(n4910) );
  OR2X1_RVT U5484 ( .A1(n12446), .A2(n4941), .Y(n5512) );
  OR2X1_RVT U5485 ( .A1(n12706), .A2(n4896), .Y(n4941) );
  OR2X1_RVT U5486 ( .A1(n5513), .A2(n4954), .Y(n5496) );
  AND4X1_RVT U5487 ( .A1(n5514), .A2(n5515), .A3(n5190), .A4(n5017), .Y(n5513)
         );
  OR2X1_RVT U5488 ( .A1(n5163), .A2(n5263), .Y(n5017) );
  OR2X1_RVT U5489 ( .A1(n4912), .A2(n5442), .Y(n5190) );
  OR2X1_RVT U5490 ( .A1(n12452), .A2(n12445), .Y(n5442) );
  OR2X1_RVT U5491 ( .A1(n296), .A2(n4834), .Y(n5515) );
  OR2X1_RVT U5492 ( .A1(n294), .A2(n12471), .Y(n5514) );
  OR2X1_RVT U5493 ( .A1(n5516), .A2(n4890), .Y(n5495) );
  AND2X1_RVT U5494 ( .A1(n5517), .A2(n4911), .Y(n5516) );
  AND2X1_RVT U5495 ( .A1(n5449), .A2(n5244), .Y(n5517) );
  OR2X1_RVT U5496 ( .A1(n5518), .A2(n12703), .Y(n5244) );
  AND2X1_RVT U5497 ( .A1(n4932), .A2(n5519), .Y(n5518) );
  OR2X1_RVT U5498 ( .A1(n12449), .A2(n4819), .Y(n5519) );
  OR2X1_RVT U5499 ( .A1(n4980), .A2(n5201), .Y(n5449) );
  OR2X1_RVT U5500 ( .A1(n4965), .A2(n4854), .Y(n5201) );
  OR2X1_RVT U5501 ( .A1(n5520), .A2(n4958), .Y(n5494) );
  AND2X1_RVT U5502 ( .A1(n5521), .A2(n12457), .Y(n5520) );
  AND2X1_RVT U5503 ( .A1(n5522), .A2(n5222), .Y(n5521) );
  OR2X1_RVT U5504 ( .A1(n4980), .A2(n5163), .Y(n5522) );
  AND4X1_RVT U5505 ( .A1(n5523), .A2(n5524), .A3(n5525), .A4(n5526), .Y(n5466)
         );
  AND2X1_RVT U5506 ( .A1(n5527), .A2(n5528), .Y(n5526) );
  OR2X1_RVT U5507 ( .A1(n12699), .A2(n5143), .Y(n5528) );
  OR2X1_RVT U5508 ( .A1(n12465), .A2(n5529), .Y(n5143) );
  OR2X1_RVT U5509 ( .A1(n4876), .A2(n4965), .Y(n5529) );
  AND2X1_RVT U5510 ( .A1(n5530), .A2(n5531), .Y(n5527) );
  OR2X1_RVT U5511 ( .A1(n4849), .A2(n4860), .Y(n5531) );
  OR2X1_RVT U5512 ( .A1(n4893), .A2(n5171), .Y(n4860) );
  OR2X1_RVT U5513 ( .A1(n12695), .A2(n4854), .Y(n5171) );
  OR2X1_RVT U5514 ( .A1(n4896), .A2(n4973), .Y(n5530) );
  OR2X1_RVT U5515 ( .A1(n4884), .A2(n5532), .Y(n4973) );
  OR2X1_RVT U5516 ( .A1(n4884), .A2(n5147), .Y(n5525) );
  OR2X1_RVT U5517 ( .A1(n296), .A2(n12467), .Y(n5147) );
  OR2X1_RVT U5518 ( .A1(n5533), .A2(n4840), .Y(n5524) );
  AND4X1_RVT U5519 ( .A1(n5534), .A2(n5535), .A3(n5536), .A4(n5537), .Y(n5533)
         );
  OR2X1_RVT U5520 ( .A1(n12693), .A2(n5538), .Y(n5536) );
  OR2X1_RVT U5521 ( .A1(n5539), .A2(n12700), .Y(n5538) );
  AND2X1_RVT U5522 ( .A1(n4891), .A2(n5540), .Y(n5539) );
  OR2X1_RVT U5523 ( .A1(n12460), .A2(n5541), .Y(n5535) );
  OR2X1_RVT U5524 ( .A1(n5280), .A2(n4834), .Y(n5541) );
  OR2X1_RVT U5525 ( .A1(n4817), .A2(n4843), .Y(n5534) );
  OR2X1_RVT U5526 ( .A1(n12697), .A2(n4943), .Y(n4843) );
  OR2X1_RVT U5527 ( .A1(n5400), .A2(n5314), .Y(n5523) );
  OR2X1_RVT U5528 ( .A1(n12476), .A2(n4854), .Y(n5314) );
  AND4X1_RVT U5529 ( .A1(n5543), .A2(n5544), .A3(n5545), .A4(n5546), .Y(n5542)
         );
  AND4X1_RVT U5530 ( .A1(n5547), .A2(n5548), .A3(n5549), .A4(n5550), .Y(n5546)
         );
  AND4X1_RVT U5531 ( .A1(n5551), .A2(n5552), .A3(n5553), .A4(n5554), .Y(n5550)
         );
  OR2X1_RVT U5532 ( .A1(n5388), .A2(n5532), .Y(n5554) );
  OR2X1_RVT U5533 ( .A1(n12696), .A2(n12470), .Y(n5532) );
  OR2X1_RVT U5534 ( .A1(n12444), .A2(n12454), .Y(n5388) );
  OR2X1_RVT U5535 ( .A1(n5555), .A2(n4891), .Y(n5553) );
  AND2X1_RVT U5536 ( .A1(n4837), .A2(n5487), .Y(n5555) );
  OR2X1_RVT U5537 ( .A1(n296), .A2(n5556), .Y(n4837) );
  OR2X1_RVT U5538 ( .A1(n12444), .A2(n12693), .Y(n5556) );
  OR2X1_RVT U5539 ( .A1(n5557), .A2(n4819), .Y(n5552) );
  OR2X1_RVT U5540 ( .A1(n12458), .A2(n4980), .Y(n4819) );
  AND2X1_RVT U5541 ( .A1(n4955), .A2(n5558), .Y(n5557) );
  OR2X1_RVT U5542 ( .A1(n4834), .A2(n5119), .Y(n5558) );
  OR2X1_RVT U5543 ( .A1(n12462), .A2(n12450), .Y(n4834) );
  OR2X1_RVT U5544 ( .A1(n5163), .A2(n5559), .Y(n4955) );
  OR2X1_RVT U5545 ( .A1(n12704), .A2(n12465), .Y(n5559) );
  OR2X1_RVT U5546 ( .A1(n5560), .A2(n4878), .Y(n5551) );
  AND2X1_RVT U5547 ( .A1(n5358), .A2(n5561), .Y(n5560) );
  OR2X1_RVT U5548 ( .A1(n5562), .A2(n12693), .Y(n5561) );
  AND2X1_RVT U5549 ( .A1(n4934), .A2(n5370), .Y(n5562) );
  OR2X1_RVT U5550 ( .A1(n12701), .A2(n4896), .Y(n5370) );
  OR2X1_RVT U5551 ( .A1(n12471), .A2(n5563), .Y(n5358) );
  OR2X1_RVT U5552 ( .A1(n12706), .A2(n12702), .Y(n5563) );
  OR2X1_RVT U5553 ( .A1(n5564), .A2(n12449), .Y(n5549) );
  AND2X1_RVT U5554 ( .A1(n5565), .A2(n5566), .Y(n5564) );
  OR2X1_RVT U5555 ( .A1(n5567), .A2(n4980), .Y(n5566) );
  AND2X1_RVT U5556 ( .A1(n5128), .A2(n5568), .Y(n5567) );
  OR2X1_RVT U5557 ( .A1(n4836), .A2(n4958), .Y(n5565) );
  OR2X1_RVT U5558 ( .A1(n12463), .A2(n4894), .Y(n4958) );
  OR2X1_RVT U5559 ( .A1(n5569), .A2(n12702), .Y(n5548) );
  AND2X1_RVT U5560 ( .A1(n5133), .A2(n5292), .Y(n5569) );
  OR2X1_RVT U5561 ( .A1(n12461), .A2(n5570), .Y(n5292) );
  OR2X1_RVT U5562 ( .A1(n4890), .A2(n12450), .Y(n5570) );
  OR2X1_RVT U5563 ( .A1(n4836), .A2(n5400), .Y(n5133) );
  OR2X1_RVT U5564 ( .A1(n12450), .A2(n12465), .Y(n5400) );
  OR2X1_RVT U5565 ( .A1(n5571), .A2(n12447), .Y(n5547) );
  AND2X1_RVT U5566 ( .A1(n5173), .A2(n5572), .Y(n5571) );
  OR2X1_RVT U5567 ( .A1(n5387), .A2(n4884), .Y(n5572) );
  OR2X1_RVT U5568 ( .A1(n4943), .A2(n5508), .Y(n5173) );
  OR2X1_RVT U5569 ( .A1(n12701), .A2(n296), .Y(n5508) );
  AND2X1_RVT U5570 ( .A1(n12451), .A2(n12704), .Y(n5269) );
  AND4X1_RVT U5571 ( .A1(n5573), .A2(n5574), .A3(n5575), .A4(n5576), .Y(n5545)
         );
  AND4X1_RVT U5572 ( .A1(n5577), .A2(n5578), .A3(n5579), .A4(n5580), .Y(n5576)
         );
  OR2X1_RVT U5573 ( .A1(n5581), .A2(n12456), .Y(n5580) );
  AND2X1_RVT U5574 ( .A1(n5160), .A2(n5231), .Y(n5581) );
  OR2X1_RVT U5575 ( .A1(n4893), .A2(n5487), .Y(n5231) );
  OR2X1_RVT U5576 ( .A1(n12704), .A2(n4890), .Y(n5487) );
  OR2X1_RVT U5577 ( .A1(n12691), .A2(n12446), .Y(n4893) );
  OR2X1_RVT U5578 ( .A1(n12447), .A2(n5263), .Y(n5160) );
  OR2X1_RVT U5579 ( .A1(n12451), .A2(n12465), .Y(n5263) );
  OR2X1_RVT U5580 ( .A1(n5582), .A2(n12700), .Y(n5579) );
  AND2X1_RVT U5581 ( .A1(n5322), .A2(n5583), .Y(n5582) );
  OR2X1_RVT U5582 ( .A1(n5280), .A2(n4907), .Y(n5583) );
  OR2X1_RVT U5583 ( .A1(n5163), .A2(n5584), .Y(n4907) );
  OR2X1_RVT U5584 ( .A1(n12476), .A2(n12452), .Y(n5584) );
  OR2X1_RVT U5585 ( .A1(n12460), .A2(n5585), .Y(n5322) );
  OR2X1_RVT U5586 ( .A1(n5163), .A2(n4876), .Y(n5585) );
  OR2X1_RVT U5587 ( .A1(n5586), .A2(n12706), .Y(n5578) );
  AND2X1_RVT U5588 ( .A1(n5268), .A2(n5197), .Y(n5586) );
  OR2X1_RVT U5589 ( .A1(n4896), .A2(n4932), .Y(n5197) );
  OR2X1_RVT U5590 ( .A1(n12698), .A2(n5163), .Y(n4932) );
  OR2X1_RVT U5591 ( .A1(n5387), .A2(n4912), .Y(n5268) );
  OR2X1_RVT U5592 ( .A1(n12457), .A2(n12703), .Y(n5387) );
  OR2X1_RVT U5593 ( .A1(n5587), .A2(n4954), .Y(n5577) );
  AND2X1_RVT U5594 ( .A1(n5588), .A2(n5589), .Y(n5587) );
  OR2X1_RVT U5595 ( .A1(n4876), .A2(n5386), .Y(n5589) );
  OR2X1_RVT U5596 ( .A1(n12700), .A2(n304), .Y(n5386) );
  AND2X1_RVT U5597 ( .A1(n5590), .A2(n5254), .Y(n5588) );
  OR2X1_RVT U5598 ( .A1(n4884), .A2(n5591), .Y(n5254) );
  OR2X1_RVT U5599 ( .A1(n12473), .A2(n12452), .Y(n5591) );
  OR2X1_RVT U5600 ( .A1(n4940), .A2(n4877), .Y(n5575) );
  OR2X1_RVT U5601 ( .A1(n12693), .A2(n4836), .Y(n4940) );
  OR2X1_RVT U5602 ( .A1(n5592), .A2(n4840), .Y(n5574) );
  AND2X1_RVT U5603 ( .A1(n5593), .A2(n5021), .Y(n5592) );
  AND2X1_RVT U5604 ( .A1(n5594), .A2(n5595), .Y(n5021) );
  OR2X1_RVT U5605 ( .A1(n12461), .A2(n5128), .Y(n5595) );
  OR2X1_RVT U5606 ( .A1(n4943), .A2(n4817), .Y(n5594) );
  OR2X1_RVT U5607 ( .A1(n12446), .A2(n4890), .Y(n4817) );
  AND2X1_RVT U5608 ( .A1(n5596), .A2(n5290), .Y(n5593) );
  OR2X1_RVT U5609 ( .A1(n4974), .A2(n5540), .Y(n5290) );
  OR2X1_RVT U5610 ( .A1(n12695), .A2(n294), .Y(n5540) );
  OR2X1_RVT U5611 ( .A1(n4836), .A2(n5003), .Y(n5596) );
  OR2X1_RVT U5612 ( .A1(n12445), .A2(n5597), .Y(n5003) );
  OR2X1_RVT U5613 ( .A1(n12691), .A2(n12474), .Y(n5597) );
  OR2X1_RVT U5614 ( .A1(n5598), .A2(n12691), .Y(n5573) );
  AND4X1_RVT U5615 ( .A1(n5599), .A2(n5600), .A3(n5601), .A4(n5432), .Y(n5598)
         );
  OR2X1_RVT U5616 ( .A1(n4890), .A2(n5353), .Y(n5432) );
  OR2X1_RVT U5617 ( .A1(n12696), .A2(n12702), .Y(n5353) );
  OR2X1_RVT U5618 ( .A1(n4890), .A2(n5602), .Y(n5601) );
  OR2X1_RVT U5619 ( .A1(n12451), .A2(n12456), .Y(n5602) );
  OR2X1_RVT U5620 ( .A1(n12701), .A2(n4849), .Y(n4890) );
  OR2X1_RVT U5621 ( .A1(n5603), .A2(n4971), .Y(n5600) );
  OR2X1_RVT U5622 ( .A1(n12445), .A2(n4815), .Y(n4971) );
  AND2X1_RVT U5623 ( .A1(n4954), .A2(n5604), .Y(n5603) );
  OR2X1_RVT U5624 ( .A1(n12699), .A2(n4854), .Y(n5604) );
  OR2X1_RVT U5625 ( .A1(n12695), .A2(n12456), .Y(n4954) );
  OR2X1_RVT U5626 ( .A1(n12697), .A2(n5568), .Y(n5599) );
  OR2X1_RVT U5627 ( .A1(n12701), .A2(n4894), .Y(n5568) );
  OR2X1_RVT U5628 ( .A1(n4840), .A2(n294), .Y(n4894) );
  AND4X1_RVT U5629 ( .A1(n5605), .A2(n5606), .A3(n5607), .A4(n5608), .Y(n5544)
         );
  AND4X1_RVT U5630 ( .A1(n5609), .A2(n5610), .A3(n5611), .A4(n5612), .Y(n5608)
         );
  OR2X1_RVT U5631 ( .A1(n4912), .A2(n5122), .Y(n5612) );
  OR2X1_RVT U5632 ( .A1(n12458), .A2(n4934), .Y(n5122) );
  OR2X1_RVT U5633 ( .A1(n12462), .A2(n5163), .Y(n4912) );
  OR2X1_RVT U5634 ( .A1(n4899), .A2(n5458), .Y(n5611) );
  OR2X1_RVT U5635 ( .A1(n12705), .A2(n12445), .Y(n5458) );
  OR2X1_RVT U5636 ( .A1(n4965), .A2(n4891), .Y(n4899) );
  OR2X1_RVT U5637 ( .A1(n4884), .A2(n4911), .Y(n5610) );
  OR2X1_RVT U5638 ( .A1(n12454), .A2(n12467), .Y(n4911) );
  OR2X1_RVT U5639 ( .A1(n12444), .A2(n12692), .Y(n4884) );
  OR2X1_RVT U5640 ( .A1(n304), .A2(n5333), .Y(n5609) );
  OR2X1_RVT U5641 ( .A1(n12452), .A2(n5120), .Y(n5333) );
  OR2X1_RVT U5642 ( .A1(n4854), .A2(n5367), .Y(n5607) );
  OR2X1_RVT U5643 ( .A1(n304), .A2(n5613), .Y(n5367) );
  OR2X1_RVT U5644 ( .A1(n12698), .A2(n12465), .Y(n5613) );
  AND2X1_RVT U5645 ( .A1(n12446), .A2(n12449), .Y(n5397) );
  OR2X1_RVT U5646 ( .A1(n4896), .A2(n4844), .Y(n5606) );
  OR2X1_RVT U5647 ( .A1(n12474), .A2(n5614), .Y(n4844) );
  OR2X1_RVT U5648 ( .A1(n12699), .A2(n12691), .Y(n5614) );
  OR2X1_RVT U5649 ( .A1(n12451), .A2(n4876), .Y(n4896) );
  OR2X1_RVT U5650 ( .A1(n4943), .A2(n5590), .Y(n5605) );
  OR2X1_RVT U5651 ( .A1(n12447), .A2(n4898), .Y(n5590) );
  OR2X1_RVT U5652 ( .A1(n12701), .A2(n12702), .Y(n4898) );
  AND4X1_RVT U5653 ( .A1(n5615), .A2(n5009), .A3(n5616), .A4(n5617), .Y(n5543)
         );
  OR2X1_RVT U5654 ( .A1(n12451), .A2(n5537), .Y(n5617) );
  OR2X1_RVT U5655 ( .A1(n12697), .A2(n5004), .Y(n5537) );
  OR2X1_RVT U5656 ( .A1(n12449), .A2(n5128), .Y(n5004) );
  OR2X1_RVT U5657 ( .A1(n12444), .A2(n4871), .Y(n5128) );
  AND2X1_RVT U5658 ( .A1(n5618), .A2(n5619), .Y(n5616) );
  OR2X1_RVT U5659 ( .A1(n12473), .A2(n5457), .Y(n5619) );
  OR2X1_RVT U5660 ( .A1(n4943), .A2(n5119), .Y(n5457) );
  OR2X1_RVT U5661 ( .A1(n12451), .A2(n12445), .Y(n5119) );
  OR2X1_RVT U5662 ( .A1(n12446), .A2(n4832), .Y(n4871) );
  OR2X1_RVT U5663 ( .A1(n12704), .A2(n5188), .Y(n5618) );
  OR2X1_RVT U5664 ( .A1(n12470), .A2(n5222), .Y(n5188) );
  OR2X1_RVT U5665 ( .A1(n12696), .A2(n12691), .Y(n5222) );
  OR2X1_RVT U5666 ( .A1(n12694), .A2(n12462), .Y(n4815) );
  AND2X1_RVT U5667 ( .A1(n5620), .A2(n5621), .Y(n5009) );
  OR2X1_RVT U5668 ( .A1(n4891), .A2(n4877), .Y(n5621) );
  OR2X1_RVT U5669 ( .A1(n12703), .A2(n4849), .Y(n4877) );
  AND2X1_RVT U5670 ( .A1(n4876), .A2(n4840), .Y(n4929) );
  OR2X1_RVT U5671 ( .A1(n12457), .A2(n4943), .Y(n4891) );
  OR2X1_RVT U5672 ( .A1(n12692), .A2(n4980), .Y(n4943) );
  OR2X1_RVT U5673 ( .A1(n5622), .A2(n4934), .Y(n5620) );
  OR2X1_RVT U5674 ( .A1(n12451), .A2(n294), .Y(n4934) );
  AND2X1_RVT U5675 ( .A1(n12705), .A2(n12444), .Y(n5280) );
  OR2X1_RVT U5676 ( .A1(n12450), .A2(n5120), .Y(n5622) );
  OR2X1_RVT U5677 ( .A1(n12701), .A2(n12467), .Y(n5120) );
  AND2X1_RVT U5678 ( .A1(n5623), .A2(n5624), .Y(n5615) );
  OR2X1_RVT U5679 ( .A1(n4857), .A2(n5273), .Y(n5624) );
  OR2X1_RVT U5680 ( .A1(n12452), .A2(n4897), .Y(n5273) );
  OR2X1_RVT U5681 ( .A1(n12467), .A2(n4974), .Y(n4897) );
  OR2X1_RVT U5682 ( .A1(n12447), .A2(n12450), .Y(n4974) );
  OR2X1_RVT U5683 ( .A1(n12698), .A2(n12696), .Y(n4836) );
  OR2X1_RVT U5684 ( .A1(n12706), .A2(n12700), .Y(n4857) );
  XOR2X1_RVT U5685 ( .A1(key[12]), .A2(state[12]), .Y(n4832) );
  OR2X1_RVT U5686 ( .A1(n4849), .A2(n4978), .Y(n5623) );
  OR2X1_RVT U5687 ( .A1(n5163), .A2(n5354), .Y(n4978) );
  OR2X1_RVT U5688 ( .A1(n12454), .A2(n4878), .Y(n5354) );
  OR2X1_RVT U5689 ( .A1(n12699), .A2(n4980), .Y(n4878) );
  XOR2X1_RVT U5690 ( .A1(key[10]), .A2(state[10]), .Y(n4980) );
  XOR2X1_RVT U5691 ( .A1(key[11]), .A2(state[11]), .Y(n4914) );
  OR2X1_RVT U5692 ( .A1(n12704), .A2(n12452), .Y(n4854) );
  XOR2X1_RVT U5693 ( .A1(key[13]), .A2(state[13]), .Y(n4840) );
  XOR2X1_RVT U5694 ( .A1(key[14]), .A2(state[14]), .Y(n4876) );
  OR2X1_RVT U5695 ( .A1(n12694), .A2(n12450), .Y(n5163) );
  XOR2X1_RVT U5696 ( .A1(key[8]), .A2(state[8]), .Y(n4855) );
  XOR2X1_RVT U5697 ( .A1(key[9]), .A2(state[9]), .Y(n4965) );
  XOR2X1_RVT U5698 ( .A1(key[15]), .A2(state[15]), .Y(n4849) );
  AND4X1_RVT U5699 ( .A1(n5626), .A2(n5627), .A3(n5628), .A4(n5629), .Y(n5625)
         );
  AND4X1_RVT U5700 ( .A1(n5630), .A2(n5631), .A3(n5632), .A4(n5633), .Y(n5629)
         );
  AND4X1_RVT U5701 ( .A1(n5634), .A2(n5635), .A3(n5636), .A4(n5637), .Y(n5633)
         );
  OR2X1_RVT U5702 ( .A1(n12438), .A2(n5639), .Y(n5632) );
  OR2X1_RVT U5703 ( .A1(n5640), .A2(n5641), .Y(n5630) );
  OR2X1_RVT U5704 ( .A1(n12688), .A2(n5642), .Y(n5641) );
  AND4X1_RVT U5705 ( .A1(n5643), .A2(n5644), .A3(n5645), .A4(n5646), .Y(n5628)
         );
  OR2X1_RVT U5706 ( .A1(n5647), .A2(n12686), .Y(n5646) );
  AND2X1_RVT U5707 ( .A1(n5648), .A2(n5649), .Y(n5647) );
  AND2X1_RVT U5708 ( .A1(n5650), .A2(n5651), .Y(n5645) );
  OR2X1_RVT U5709 ( .A1(n5652), .A2(n316), .Y(n5651) );
  AND2X1_RVT U5710 ( .A1(n5653), .A2(n5654), .Y(n5652) );
  OR2X1_RVT U5711 ( .A1(n12429), .A2(n5656), .Y(n5654) );
  OR2X1_RVT U5712 ( .A1(n5642), .A2(n5657), .Y(n5653) );
  OR2X1_RVT U5713 ( .A1(n5658), .A2(n12435), .Y(n5650) );
  AND2X1_RVT U5714 ( .A1(n5660), .A2(n5661), .Y(n5658) );
  OR2X1_RVT U5715 ( .A1(n5662), .A2(n5663), .Y(n5644) );
  AND2X1_RVT U5716 ( .A1(n5664), .A2(n5665), .Y(n5662) );
  OR2X1_RVT U5717 ( .A1(n12430), .A2(n5666), .Y(n5665) );
  AND2X1_RVT U5718 ( .A1(n5667), .A2(n5668), .Y(n5664) );
  AND2X1_RVT U5719 ( .A1(n5669), .A2(n5670), .Y(n5643) );
  OR2X1_RVT U5720 ( .A1(n5671), .A2(n12412), .Y(n5670) );
  AND2X1_RVT U5721 ( .A1(n5673), .A2(n5674), .Y(n5671) );
  OR2X1_RVT U5722 ( .A1(n5675), .A2(n5676), .Y(n5674) );
  OR2X1_RVT U5723 ( .A1(n12421), .A2(n12416), .Y(n5676) );
  OR2X1_RVT U5724 ( .A1(n5679), .A2(n5680), .Y(n5669) );
  AND2X1_RVT U5725 ( .A1(n5681), .A2(n5682), .Y(n5679) );
  AND2X1_RVT U5726 ( .A1(n5683), .A2(n5684), .Y(n5681) );
  AND4X1_RVT U5727 ( .A1(n5685), .A2(n5686), .A3(n5687), .A4(n5688), .Y(n5627)
         );
  AND4X1_RVT U5728 ( .A1(n5689), .A2(n5690), .A3(n5691), .A4(n5692), .Y(n5688)
         );
  OR2X1_RVT U5729 ( .A1(n5693), .A2(n12441), .Y(n5692) );
  AND4X1_RVT U5730 ( .A1(n5695), .A2(n5696), .A3(n5697), .A4(n5698), .Y(n5693)
         );
  OR2X1_RVT U5731 ( .A1(n5699), .A2(n5666), .Y(n5698) );
  OR2X1_RVT U5732 ( .A1(n5700), .A2(n12427), .Y(n5697) );
  OR2X1_RVT U5733 ( .A1(n5702), .A2(n12418), .Y(n5691) );
  AND4X1_RVT U5734 ( .A1(n5703), .A2(n5704), .A3(n5705), .A4(n5706), .Y(n5702)
         );
  OR2X1_RVT U5735 ( .A1(n5707), .A2(n5708), .Y(n5706) );
  OR2X1_RVT U5736 ( .A1(n12435), .A2(n12430), .Y(n5708) );
  AND2X1_RVT U5737 ( .A1(n5709), .A2(n5710), .Y(n5705) );
  OR2X1_RVT U5738 ( .A1(n12690), .A2(n5711), .Y(n5704) );
  OR2X1_RVT U5739 ( .A1(n5712), .A2(n5713), .Y(n5703) );
  AND2X1_RVT U5740 ( .A1(n5714), .A2(n5715), .Y(n5712) );
  OR2X1_RVT U5741 ( .A1(n12435), .A2(n5716), .Y(n5715) );
  OR2X1_RVT U5742 ( .A1(n5649), .A2(n5717), .Y(n5690) );
  OR2X1_RVT U5743 ( .A1(n5716), .A2(n5718), .Y(n5689) );
  OR2X1_RVT U5744 ( .A1(n5719), .A2(n5720), .Y(n5687) );
  OR2X1_RVT U5745 ( .A1(n5721), .A2(n5714), .Y(n5686) );
  OR2X1_RVT U5746 ( .A1(n5722), .A2(n5723), .Y(n5685) );
  AND4X1_RVT U5747 ( .A1(n5724), .A2(n5725), .A3(n5726), .A4(n5727), .Y(n5626)
         );
  AND2X1_RVT U5748 ( .A1(n5728), .A2(n5729), .Y(n5727) );
  OR2X1_RVT U5749 ( .A1(n5713), .A2(n5730), .Y(n5729) );
  AND2X1_RVT U5750 ( .A1(n5731), .A2(n5732), .Y(n5728) );
  OR2X1_RVT U5751 ( .A1(n5733), .A2(n5656), .Y(n5732) );
  OR2X1_RVT U5752 ( .A1(n5657), .A2(n5734), .Y(n5731) );
  OR2X1_RVT U5753 ( .A1(n314), .A2(n5735), .Y(n5726) );
  OR2X1_RVT U5754 ( .A1(n5736), .A2(n12425), .Y(n5725) );
  OR2X1_RVT U5755 ( .A1(n12428), .A2(n5738), .Y(n5724) );
  AND4X1_RVT U5756 ( .A1(n5740), .A2(n5741), .A3(n5742), .A4(n5743), .Y(n5739)
         );
  AND4X1_RVT U5757 ( .A1(n5744), .A2(n5635), .A3(n5745), .A4(n5746), .Y(n5743)
         );
  AND4X1_RVT U5758 ( .A1(n5747), .A2(n5748), .A3(n5749), .A4(n5750), .Y(n5746)
         );
  OR2X1_RVT U5759 ( .A1(n5656), .A2(n5751), .Y(n5750) );
  OR2X1_RVT U5760 ( .A1(n5752), .A2(n12440), .Y(n5751) );
  OR2X1_RVT U5761 ( .A1(n5657), .A2(n5753), .Y(n5749) );
  OR2X1_RVT U5762 ( .A1(n314), .A2(n12424), .Y(n5753) );
  OR2X1_RVT U5763 ( .A1(n5754), .A2(n5700), .Y(n5748) );
  AND2X1_RVT U5764 ( .A1(n5711), .A2(n5755), .Y(n5754) );
  OR2X1_RVT U5765 ( .A1(n5756), .A2(n5757), .Y(n5747) );
  AND2X1_RVT U5766 ( .A1(n5758), .A2(n5759), .Y(n5756) );
  AND2X1_RVT U5767 ( .A1(n5760), .A2(n5761), .Y(n5745) );
  OR2X1_RVT U5768 ( .A1(n5707), .A2(n5762), .Y(n5761) );
  OR2X1_RVT U5769 ( .A1(n5763), .A2(n12688), .Y(n5762) );
  OR2X1_RVT U5770 ( .A1(n5764), .A2(n5765), .Y(n5760) );
  OR2X1_RVT U5771 ( .A1(n5766), .A2(n12429), .Y(n5765) );
  OR2X1_RVT U5772 ( .A1(n5642), .A2(n5767), .Y(n5635) );
  AND4X1_RVT U5773 ( .A1(n5768), .A2(n5769), .A3(n5770), .A4(n5771), .Y(n5742)
         );
  AND4X1_RVT U5774 ( .A1(n5772), .A2(n5773), .A3(n5774), .A4(n5775), .Y(n5771)
         );
  OR2X1_RVT U5775 ( .A1(n5776), .A2(n12443), .Y(n5775) );
  AND2X1_RVT U5776 ( .A1(n5778), .A2(n5779), .Y(n5776) );
  OR2X1_RVT U5777 ( .A1(n12412), .A2(n5657), .Y(n5779) );
  OR2X1_RVT U5778 ( .A1(n5780), .A2(n5659), .Y(n5774) );
  AND2X1_RVT U5779 ( .A1(n5781), .A2(n5782), .Y(n5780) );
  OR2X1_RVT U5780 ( .A1(n5783), .A2(n12687), .Y(n5773) );
  AND2X1_RVT U5781 ( .A1(n5784), .A2(n5785), .Y(n5783) );
  OR2X1_RVT U5782 ( .A1(n5786), .A2(n5735), .Y(n5785) );
  AND2X1_RVT U5783 ( .A1(n12443), .A2(n12427), .Y(n5786) );
  OR2X1_RVT U5784 ( .A1(n5787), .A2(n12413), .Y(n5772) );
  AND2X1_RVT U5785 ( .A1(n5789), .A2(n5790), .Y(n5787) );
  OR2X1_RVT U5786 ( .A1(n5791), .A2(n12419), .Y(n5770) );
  AND2X1_RVT U5787 ( .A1(n5792), .A2(n5793), .Y(n5791) );
  OR2X1_RVT U5788 ( .A1(n12427), .A2(n5794), .Y(n5793) );
  AND2X1_RVT U5789 ( .A1(n5795), .A2(n5796), .Y(n5792) );
  OR2X1_RVT U5790 ( .A1(n5797), .A2(n5798), .Y(n5795) );
  OR2X1_RVT U5791 ( .A1(n5642), .A2(n5713), .Y(n5798) );
  OR2X1_RVT U5792 ( .A1(n5799), .A2(n12684), .Y(n5769) );
  AND2X1_RVT U5793 ( .A1(n5800), .A2(n5801), .Y(n5799) );
  OR2X1_RVT U5794 ( .A1(n5802), .A2(n5803), .Y(n5768) );
  AND2X1_RVT U5795 ( .A1(n5804), .A2(n5805), .Y(n5802) );
  AND2X1_RVT U5796 ( .A1(n5806), .A2(n5807), .Y(n5804) );
  OR2X1_RVT U5797 ( .A1(n316), .A2(n5735), .Y(n5807) );
  OR2X1_RVT U5798 ( .A1(n12437), .A2(n5700), .Y(n5806) );
  AND4X1_RVT U5799 ( .A1(n5808), .A2(n5809), .A3(n5810), .A4(n5811), .Y(n5741)
         );
  AND4X1_RVT U5800 ( .A1(n5812), .A2(n5813), .A3(n5814), .A4(n5815), .Y(n5811)
         );
  OR2X1_RVT U5801 ( .A1(n5735), .A2(n5734), .Y(n5815) );
  OR2X1_RVT U5802 ( .A1(n5666), .A2(n5816), .Y(n5814) );
  OR2X1_RVT U5803 ( .A1(n5699), .A2(n5817), .Y(n5813) );
  OR2X1_RVT U5804 ( .A1(n5642), .A2(n5818), .Y(n5812) );
  AND2X1_RVT U5805 ( .A1(n5819), .A2(n5820), .Y(n5810) );
  OR2X1_RVT U5806 ( .A1(n12438), .A2(n5821), .Y(n5820) );
  OR2X1_RVT U5807 ( .A1(n12417), .A2(n5718), .Y(n5819) );
  OR2X1_RVT U5808 ( .A1(n5822), .A2(n5677), .Y(n5809) );
  AND4X1_RVT U5809 ( .A1(n5823), .A2(n5824), .A3(n5825), .A4(n5826), .Y(n5822)
         );
  OR2X1_RVT U5810 ( .A1(n5827), .A2(n5642), .Y(n5825) );
  OR2X1_RVT U5811 ( .A1(n12676), .A2(n5828), .Y(n5824) );
  OR2X1_RVT U5812 ( .A1(n5829), .A2(n12684), .Y(n5823) );
  AND2X1_RVT U5813 ( .A1(n5720), .A2(n5830), .Y(n5829) );
  OR2X1_RVT U5814 ( .A1(n5722), .A2(n5831), .Y(n5808) );
  AND4X1_RVT U5815 ( .A1(n5832), .A2(n5833), .A3(n5834), .A4(n5835), .Y(n5740)
         );
  AND4X1_RVT U5816 ( .A1(n5836), .A2(n5837), .A3(n5838), .A4(n5839), .Y(n5835)
         );
  OR2X1_RVT U5817 ( .A1(n12680), .A2(n5840), .Y(n5839) );
  OR2X1_RVT U5818 ( .A1(n12681), .A2(n5841), .Y(n5838) );
  OR2X1_RVT U5819 ( .A1(n12678), .A2(n5842), .Y(n5837) );
  OR2X1_RVT U5820 ( .A1(n12411), .A2(n5843), .Y(n5836) );
  OR2X1_RVT U5821 ( .A1(n5844), .A2(n12418), .Y(n5833) );
  AND4X1_RVT U5822 ( .A1(n5846), .A2(n5847), .A3(n5848), .A4(n5849), .Y(n5845)
         );
  AND4X1_RVT U5823 ( .A1(n5850), .A2(n5851), .A3(n5852), .A4(n5853), .Y(n5849)
         );
  AND4X1_RVT U5824 ( .A1(n5854), .A2(n5631), .A3(n5801), .A4(n5855), .Y(n5853)
         );
  OR2X1_RVT U5825 ( .A1(n5856), .A2(n12675), .Y(n5631) );
  AND2X1_RVT U5826 ( .A1(n5857), .A2(n5858), .Y(n5856) );
  OR2X1_RVT U5827 ( .A1(n5675), .A2(n5859), .Y(n5858) );
  OR2X1_RVT U5828 ( .A1(n5860), .A2(n5757), .Y(n5857) );
  OR2X1_RVT U5829 ( .A1(n5861), .A2(n5716), .Y(n5854) );
  AND2X1_RVT U5830 ( .A1(n5862), .A2(n5863), .Y(n5861) );
  OR2X1_RVT U5831 ( .A1(n12680), .A2(n5700), .Y(n5863) );
  OR2X1_RVT U5832 ( .A1(n5864), .A2(n5659), .Y(n5852) );
  AND2X1_RVT U5833 ( .A1(n5865), .A2(n5866), .Y(n5864) );
  OR2X1_RVT U5834 ( .A1(n5867), .A2(n12686), .Y(n5866) );
  AND2X1_RVT U5835 ( .A1(n5707), .A2(n5868), .Y(n5867) );
  OR2X1_RVT U5836 ( .A1(n5869), .A2(n12438), .Y(n5851) );
  AND2X1_RVT U5837 ( .A1(n5870), .A2(n5871), .Y(n5869) );
  OR2X1_RVT U5838 ( .A1(n5700), .A2(n5666), .Y(n5871) );
  OR2X1_RVT U5839 ( .A1(n5872), .A2(n12421), .Y(n5850) );
  AND2X1_RVT U5840 ( .A1(n5784), .A2(n5873), .Y(n5872) );
  OR2X1_RVT U5841 ( .A1(n5713), .A2(n5874), .Y(n5784) );
  AND4X1_RVT U5842 ( .A1(n5875), .A2(n5876), .A3(n5877), .A4(n5878), .Y(n5848)
         );
  OR2X1_RVT U5843 ( .A1(n5879), .A2(n12428), .Y(n5878) );
  AND2X1_RVT U5844 ( .A1(n5880), .A2(n5881), .Y(n5879) );
  OR2X1_RVT U5845 ( .A1(n5757), .A2(n5657), .Y(n5881) );
  AND2X1_RVT U5846 ( .A1(n5882), .A2(n5883), .Y(n5880) );
  OR2X1_RVT U5847 ( .A1(n5797), .A2(n5859), .Y(n5882) );
  AND2X1_RVT U5848 ( .A1(n5884), .A2(n5885), .Y(n5877) );
  OR2X1_RVT U5849 ( .A1(n5886), .A2(n5788), .Y(n5885) );
  AND2X1_RVT U5850 ( .A1(n5887), .A2(n5696), .Y(n5886) );
  OR2X1_RVT U5851 ( .A1(n5642), .A2(n5757), .Y(n5696) );
  OR2X1_RVT U5852 ( .A1(n5888), .A2(n316), .Y(n5884) );
  AND2X1_RVT U5853 ( .A1(n5889), .A2(n5890), .Y(n5888) );
  OR2X1_RVT U5854 ( .A1(n5891), .A2(n12430), .Y(n5890) );
  AND2X1_RVT U5855 ( .A1(n5892), .A2(n5893), .Y(n5891) );
  OR2X1_RVT U5856 ( .A1(n12425), .A2(n5707), .Y(n5893) );
  OR2X1_RVT U5857 ( .A1(n12690), .A2(n12427), .Y(n5892) );
  AND2X1_RVT U5858 ( .A1(n5758), .A2(n5868), .Y(n5889) );
  OR2X1_RVT U5859 ( .A1(n5788), .A2(n5894), .Y(n5758) );
  OR2X1_RVT U5860 ( .A1(n12685), .A2(n12681), .Y(n5894) );
  OR2X1_RVT U5861 ( .A1(n5895), .A2(n5777), .Y(n5876) );
  AND4X1_RVT U5862 ( .A1(n5736), .A2(n5896), .A3(n5897), .A4(n5898), .Y(n5895)
         );
  OR2X1_RVT U5863 ( .A1(n12429), .A2(n5757), .Y(n5898) );
  AND2X1_RVT U5864 ( .A1(n5899), .A2(n5900), .Y(n5897) );
  OR2X1_RVT U5865 ( .A1(n12690), .A2(n12438), .Y(n5896) );
  AND2X1_RVT U5866 ( .A1(n5901), .A2(n5902), .Y(n5736) );
  OR2X1_RVT U5867 ( .A1(n5903), .A2(n314), .Y(n5902) );
  OR2X1_RVT U5868 ( .A1(n5700), .A2(n12675), .Y(n5901) );
  AND2X1_RVT U5869 ( .A1(n5904), .A2(n5905), .Y(n5875) );
  OR2X1_RVT U5870 ( .A1(n5906), .A2(n12677), .Y(n5905) );
  AND2X1_RVT U5871 ( .A1(n5907), .A2(n5908), .Y(n5906) );
  OR2X1_RVT U5872 ( .A1(n5909), .A2(n12432), .Y(n5908) );
  AND2X1_RVT U5873 ( .A1(n5910), .A2(n5911), .Y(n5909) );
  AND2X1_RVT U5874 ( .A1(n5912), .A2(n5913), .Y(n5907) );
  OR2X1_RVT U5875 ( .A1(n5914), .A2(n12441), .Y(n5904) );
  AND4X1_RVT U5876 ( .A1(n5915), .A2(n5916), .A3(n5917), .A4(n5918), .Y(n5914)
         );
  OR2X1_RVT U5877 ( .A1(n12689), .A2(n5919), .Y(n5917) );
  OR2X1_RVT U5878 ( .A1(n314), .A2(n5714), .Y(n5916) );
  OR2X1_RVT U5879 ( .A1(n5803), .A2(n5757), .Y(n5915) );
  AND4X1_RVT U5880 ( .A1(n5920), .A2(n5921), .A3(n5922), .A4(n5923), .Y(n5847)
         );
  AND2X1_RVT U5881 ( .A1(n5924), .A2(n5767), .Y(n5923) );
  OR2X1_RVT U5882 ( .A1(n12416), .A2(n5733), .Y(n5767) );
  AND2X1_RVT U5883 ( .A1(n5925), .A2(n5926), .Y(n5924) );
  OR2X1_RVT U5884 ( .A1(n5927), .A2(n5682), .Y(n5926) );
  OR2X1_RVT U5885 ( .A1(n5734), .A2(n5794), .Y(n5925) );
  OR2X1_RVT U5886 ( .A1(n314), .A2(n5928), .Y(n5922) );
  OR2X1_RVT U5887 ( .A1(n12688), .A2(n5929), .Y(n5921) );
  OR2X1_RVT U5888 ( .A1(n5803), .A2(n5930), .Y(n5920) );
  AND4X1_RVT U5889 ( .A1(n5931), .A2(n5932), .A3(n5933), .A4(n5934), .Y(n5846)
         );
  AND2X1_RVT U5890 ( .A1(n5935), .A2(n5936), .Y(n5934) );
  OR2X1_RVT U5891 ( .A1(n12411), .A2(n5937), .Y(n5936) );
  AND2X1_RVT U5892 ( .A1(n5938), .A2(n5939), .Y(n5935) );
  OR2X1_RVT U5893 ( .A1(n5699), .A2(n5709), .Y(n5939) );
  OR2X1_RVT U5894 ( .A1(n12432), .A2(n5759), .Y(n5709) );
  OR2X1_RVT U5895 ( .A1(n12418), .A2(n5940), .Y(n5938) );
  OR2X1_RVT U5896 ( .A1(n5680), .A2(n5673), .Y(n5933) );
  OR2X1_RVT U5897 ( .A1(n5766), .A2(n5941), .Y(n5673) );
  OR2X1_RVT U5898 ( .A1(n12684), .A2(n5942), .Y(n5932) );
  OR2X1_RVT U5899 ( .A1(n12430), .A2(n5800), .Y(n5931) );
  OR2X1_RVT U5900 ( .A1(n12675), .A2(n5862), .Y(n5800) );
  AND4X1_RVT U5901 ( .A1(n5944), .A2(n5945), .A3(n5946), .A4(n5947), .Y(n5943)
         );
  AND4X1_RVT U5902 ( .A1(n5948), .A2(n5949), .A3(n5950), .A4(n5951), .Y(n5947)
         );
  OR2X1_RVT U5903 ( .A1(n324), .A2(n5952), .Y(n5951) );
  OR2X1_RVT U5904 ( .A1(n5953), .A2(n12443), .Y(n5952) );
  AND2X1_RVT U5905 ( .A1(n12432), .A2(n5719), .Y(n5953) );
  AND2X1_RVT U5906 ( .A1(n5634), .A2(n5954), .Y(n5950) );
  OR2X1_RVT U5907 ( .A1(n12421), .A2(n5955), .Y(n5634) );
  OR2X1_RVT U5908 ( .A1(n324), .A2(n5713), .Y(n5955) );
  OR2X1_RVT U5909 ( .A1(n5956), .A2(n5642), .Y(n5949) );
  AND2X1_RVT U5910 ( .A1(n5957), .A2(n5958), .Y(n5956) );
  AND2X1_RVT U5911 ( .A1(n5959), .A2(n5960), .Y(n5948) );
  OR2X1_RVT U5912 ( .A1(n5961), .A2(n5962), .Y(n5960) );
  AND2X1_RVT U5913 ( .A1(n5963), .A2(n5723), .Y(n5961) );
  OR2X1_RVT U5914 ( .A1(n5964), .A2(n5714), .Y(n5959) );
  AND2X1_RVT U5915 ( .A1(n5899), .A2(n5733), .Y(n5964) );
  OR2X1_RVT U5916 ( .A1(n12419), .A2(n5965), .Y(n5899) );
  OR2X1_RVT U5917 ( .A1(n12690), .A2(n12429), .Y(n5965) );
  AND4X1_RVT U5918 ( .A1(n5966), .A2(n5967), .A3(n5968), .A4(n5969), .Y(n5946)
         );
  OR2X1_RVT U5919 ( .A1(n5970), .A2(n12680), .Y(n5969) );
  AND2X1_RVT U5920 ( .A1(n5782), .A2(n5971), .Y(n5970) );
  OR2X1_RVT U5921 ( .A1(n12688), .A2(n5827), .Y(n5782) );
  AND2X1_RVT U5922 ( .A1(n5972), .A2(n5973), .Y(n5968) );
  OR2X1_RVT U5923 ( .A1(n5974), .A2(n12678), .Y(n5973) );
  AND2X1_RVT U5924 ( .A1(n5975), .A2(n5976), .Y(n5974) );
  OR2X1_RVT U5925 ( .A1(n5677), .A2(n5919), .Y(n5976) );
  OR2X1_RVT U5926 ( .A1(n5977), .A2(n12676), .Y(n5972) );
  AND2X1_RVT U5927 ( .A1(n5978), .A2(n5979), .Y(n5977) );
  OR2X1_RVT U5928 ( .A1(n5980), .A2(n12432), .Y(n5967) );
  AND2X1_RVT U5929 ( .A1(n5981), .A2(n5982), .Y(n5980) );
  AND2X1_RVT U5930 ( .A1(n5983), .A2(n5984), .Y(n5981) );
  AND2X1_RVT U5931 ( .A1(n5985), .A2(n5986), .Y(n5966) );
  OR2X1_RVT U5932 ( .A1(n5987), .A2(n5903), .Y(n5986) );
  AND2X1_RVT U5933 ( .A1(n5988), .A2(n5734), .Y(n5987) );
  AND2X1_RVT U5934 ( .A1(n5989), .A2(n5990), .Y(n5988) );
  OR2X1_RVT U5935 ( .A1(n5991), .A2(n12435), .Y(n5985) );
  AND2X1_RVT U5936 ( .A1(n5992), .A2(n5993), .Y(n5991) );
  OR2X1_RVT U5937 ( .A1(n12687), .A2(n12437), .Y(n5993) );
  AND2X1_RVT U5938 ( .A1(n5723), .A2(n5994), .Y(n5992) );
  AND4X1_RVT U5939 ( .A1(n5995), .A2(n5996), .A3(n5997), .A4(n5998), .Y(n5945)
         );
  AND2X1_RVT U5940 ( .A1(n5999), .A2(n6000), .Y(n5998) );
  OR2X1_RVT U5941 ( .A1(n5716), .A2(n5790), .Y(n6000) );
  OR2X1_RVT U5942 ( .A1(n12682), .A2(n5723), .Y(n5790) );
  AND2X1_RVT U5943 ( .A1(n6001), .A2(n6002), .Y(n5999) );
  OR2X1_RVT U5944 ( .A1(n5868), .A2(n5682), .Y(n6002) );
  OR2X1_RVT U5945 ( .A1(n12689), .A2(n12428), .Y(n5682) );
  OR2X1_RVT U5946 ( .A1(n5766), .A2(n5816), .Y(n6001) );
  OR2X1_RVT U5947 ( .A1(n12677), .A2(n6003), .Y(n5816) );
  OR2X1_RVT U5948 ( .A1(n6004), .A2(n12411), .Y(n5997) );
  AND4X1_RVT U5949 ( .A1(n6005), .A2(n6006), .A3(n6007), .A4(n6008), .Y(n6004)
         );
  OR2X1_RVT U5950 ( .A1(n5941), .A2(n5714), .Y(n6007) );
  OR2X1_RVT U5951 ( .A1(n6009), .A2(n5711), .Y(n6006) );
  OR2X1_RVT U5952 ( .A1(n12686), .A2(n5666), .Y(n6005) );
  OR2X1_RVT U5953 ( .A1(n6010), .A2(n12412), .Y(n5996) );
  AND2X1_RVT U5954 ( .A1(n6011), .A2(n6012), .Y(n6010) );
  OR2X1_RVT U5955 ( .A1(n5941), .A2(n5666), .Y(n6012) );
  AND2X1_RVT U5956 ( .A1(n6013), .A2(n5942), .Y(n6011) );
  OR2X1_RVT U5957 ( .A1(n5714), .A2(n6014), .Y(n5942) );
  OR2X1_RVT U5958 ( .A1(n12677), .A2(n12689), .Y(n6014) );
  OR2X1_RVT U5959 ( .A1(n6015), .A2(n12419), .Y(n5995) );
  AND4X1_RVT U5960 ( .A1(n6016), .A2(n5929), .A3(n5738), .A4(n5710), .Y(n6015)
         );
  OR2X1_RVT U5961 ( .A1(n5735), .A2(n6017), .Y(n5710) );
  OR2X1_RVT U5962 ( .A1(n12679), .A2(n5672), .Y(n6017) );
  OR2X1_RVT U5963 ( .A1(n5797), .A2(n5831), .Y(n5738) );
  OR2X1_RVT U5964 ( .A1(n5716), .A2(n6018), .Y(n5929) );
  OR2X1_RVT U5965 ( .A1(n12443), .A2(n12412), .Y(n6018) );
  OR2X1_RVT U5966 ( .A1(n5675), .A2(n6019), .Y(n6016) );
  OR2X1_RVT U5967 ( .A1(n6020), .A2(n12417), .Y(n6019) );
  AND4X1_RVT U5968 ( .A1(n6021), .A2(n6022), .A3(n6023), .A4(n6024), .Y(n5944)
         );
  AND2X1_RVT U5969 ( .A1(n6025), .A2(n6026), .Y(n6024) );
  AND2X1_RVT U5970 ( .A1(n6027), .A2(n6028), .Y(n6025) );
  OR2X1_RVT U5971 ( .A1(n5707), .A2(n5982), .Y(n6028) );
  OR2X1_RVT U5972 ( .A1(n5719), .A2(n6029), .Y(n5982) );
  OR2X1_RVT U5973 ( .A1(n12678), .A2(n12680), .Y(n6029) );
  OR2X1_RVT U5974 ( .A1(n12685), .A2(n6030), .Y(n6027) );
  OR2X1_RVT U5975 ( .A1(n12428), .A2(n6031), .Y(n6023) );
  OR2X1_RVT U5976 ( .A1(n12688), .A2(n6032), .Y(n6022) );
  OR2X1_RVT U5977 ( .A1(n5719), .A2(n6033), .Y(n6021) );
  AND4X1_RVT U5978 ( .A1(n6035), .A2(n6036), .A3(n6037), .A4(n6038), .Y(n6034)
         );
  AND4X1_RVT U5979 ( .A1(n6039), .A2(n6040), .A3(n6041), .A4(n6042), .Y(n6038)
         );
  AND4X1_RVT U5980 ( .A1(n6043), .A2(n6044), .A3(n5636), .A4(n6045), .Y(n6042)
         );
  OR2X1_RVT U5981 ( .A1(n5777), .A2(n6046), .Y(n5636) );
  OR2X1_RVT U5982 ( .A1(n5868), .A2(n316), .Y(n6046) );
  OR2X1_RVT U5983 ( .A1(n5640), .A2(n6047), .Y(n6044) );
  OR2X1_RVT U5984 ( .A1(n12683), .A2(n12686), .Y(n6047) );
  OR2X1_RVT U5985 ( .A1(n5903), .A2(n6048), .Y(n6043) );
  OR2X1_RVT U5986 ( .A1(n6049), .A2(n5677), .Y(n6048) );
  AND2X1_RVT U5987 ( .A1(n12432), .A2(n5777), .Y(n6049) );
  OR2X1_RVT U5988 ( .A1(n6050), .A2(n12438), .Y(n6041) );
  AND2X1_RVT U5989 ( .A1(n5918), .A2(n5990), .Y(n6050) );
  OR2X1_RVT U5990 ( .A1(n316), .A2(n6051), .Y(n5990) );
  OR2X1_RVT U5991 ( .A1(n12411), .A2(n12682), .Y(n6051) );
  OR2X1_RVT U5992 ( .A1(n5707), .A2(n6052), .Y(n5918) );
  OR2X1_RVT U5993 ( .A1(n12680), .A2(n5699), .Y(n6052) );
  OR2X1_RVT U5994 ( .A1(n6053), .A2(n5657), .Y(n6040) );
  AND2X1_RVT U5995 ( .A1(n6054), .A2(n5862), .Y(n6053) );
  OR2X1_RVT U5996 ( .A1(n5763), .A2(n5757), .Y(n6039) );
  AND4X1_RVT U5997 ( .A1(n6055), .A2(n6056), .A3(n6057), .A4(n6058), .Y(n6037)
         );
  AND2X1_RVT U5998 ( .A1(n6059), .A2(n6060), .Y(n6058) );
  OR2X1_RVT U5999 ( .A1(n6061), .A2(n12432), .Y(n6060) );
  AND2X1_RVT U6000 ( .A1(n6062), .A2(n5730), .Y(n6061) );
  AND2X1_RVT U6001 ( .A1(n6063), .A2(n6064), .Y(n6059) );
  OR2X1_RVT U6002 ( .A1(n6065), .A2(n5713), .Y(n6064) );
  AND2X1_RVT U6003 ( .A1(n5684), .A2(n5656), .Y(n6065) );
  OR2X1_RVT U6004 ( .A1(n12688), .A2(n5755), .Y(n5684) );
  OR2X1_RVT U6005 ( .A1(n6066), .A2(n5766), .Y(n6063) );
  AND2X1_RVT U6006 ( .A1(n5958), .A2(n6067), .Y(n6066) );
  OR2X1_RVT U6007 ( .A1(n12689), .A2(n5794), .Y(n5958) );
  OR2X1_RVT U6008 ( .A1(n6068), .A2(n12680), .Y(n6057) );
  AND2X1_RVT U6009 ( .A1(n5661), .A2(n6069), .Y(n6068) );
  OR2X1_RVT U6010 ( .A1(n5797), .A2(n5721), .Y(n6069) );
  OR2X1_RVT U6011 ( .A1(n5700), .A2(n5903), .Y(n5661) );
  OR2X1_RVT U6012 ( .A1(n6070), .A2(n314), .Y(n6056) );
  AND2X1_RVT U6013 ( .A1(n5711), .A2(n6071), .Y(n6070) );
  OR2X1_RVT U6014 ( .A1(n6072), .A2(n12416), .Y(n6071) );
  AND2X1_RVT U6015 ( .A1(n6073), .A2(n6074), .Y(n6072) );
  OR2X1_RVT U6016 ( .A1(n12681), .A2(n5694), .Y(n6074) );
  OR2X1_RVT U6017 ( .A1(n12443), .A2(n5797), .Y(n5711) );
  OR2X1_RVT U6018 ( .A1(n6075), .A2(n5781), .Y(n6055) );
  AND2X1_RVT U6019 ( .A1(n5714), .A2(n5759), .Y(n6075) );
  OR2X1_RVT U6020 ( .A1(n12677), .A2(n5642), .Y(n5759) );
  AND4X1_RVT U6021 ( .A1(n6076), .A2(n6077), .A3(n6078), .A4(n6079), .Y(n6036)
         );
  AND4X1_RVT U6022 ( .A1(n6080), .A2(n6081), .A3(n6082), .A4(n6083), .Y(n6079)
         );
  OR2X1_RVT U6023 ( .A1(n6084), .A2(n12688), .Y(n6083) );
  AND2X1_RVT U6024 ( .A1(n5817), .A2(n6085), .Y(n6084) );
  OR2X1_RVT U6025 ( .A1(n12440), .A2(n5666), .Y(n6085) );
  OR2X1_RVT U6026 ( .A1(n6086), .A2(n5659), .Y(n6082) );
  AND2X1_RVT U6027 ( .A1(n6087), .A2(n6088), .Y(n6086) );
  OR2X1_RVT U6028 ( .A1(n6089), .A2(n5694), .Y(n6088) );
  AND2X1_RVT U6029 ( .A1(n5719), .A2(n5707), .Y(n6089) );
  AND2X1_RVT U6030 ( .A1(n5721), .A2(n5963), .Y(n6087) );
  OR2X1_RVT U6031 ( .A1(n12441), .A2(n5859), .Y(n5963) );
  OR2X1_RVT U6032 ( .A1(n6090), .A2(n12430), .Y(n6081) );
  AND2X1_RVT U6033 ( .A1(n6091), .A2(n6092), .Y(n6090) );
  OR2X1_RVT U6034 ( .A1(n5707), .A2(n6093), .Y(n6092) );
  AND2X1_RVT U6035 ( .A1(n5789), .A2(n5983), .Y(n6091) );
  OR2X1_RVT U6036 ( .A1(n5699), .A2(n5874), .Y(n5983) );
  OR2X1_RVT U6037 ( .A1(n5672), .A2(n6094), .Y(n5789) );
  OR2X1_RVT U6038 ( .A1(n6095), .A2(n5642), .Y(n6080) );
  AND4X1_RVT U6039 ( .A1(n6096), .A2(n6097), .A3(n6098), .A4(n6031), .Y(n6095)
         );
  OR2X1_RVT U6040 ( .A1(n5735), .A2(n6099), .Y(n6031) );
  OR2X1_RVT U6041 ( .A1(n12411), .A2(n5699), .Y(n6099) );
  OR2X1_RVT U6042 ( .A1(n12685), .A2(n5941), .Y(n6097) );
  OR2X1_RVT U6043 ( .A1(n5700), .A2(n5797), .Y(n6096) );
  OR2X1_RVT U6044 ( .A1(n5868), .A2(n5910), .Y(n6078) );
  OR2X1_RVT U6045 ( .A1(n6100), .A2(n12414), .Y(n6077) );
  AND4X1_RVT U6046 ( .A1(n6101), .A2(n6102), .A3(n5744), .A4(n5842), .Y(n6100)
         );
  OR2X1_RVT U6047 ( .A1(n5666), .A2(n5831), .Y(n5842) );
  OR2X1_RVT U6048 ( .A1(n12685), .A2(n314), .Y(n5831) );
  OR2X1_RVT U6049 ( .A1(n5659), .A2(n5723), .Y(n5744) );
  OR2X1_RVT U6050 ( .A1(n12677), .A2(n6094), .Y(n6076) );
  AND4X1_RVT U6051 ( .A1(n6103), .A2(n6104), .A3(n6105), .A4(n6106), .Y(n6035)
         );
  OR2X1_RVT U6052 ( .A1(n12419), .A2(n6107), .Y(n6106) );
  AND2X1_RVT U6053 ( .A1(n6108), .A2(n6109), .Y(n6105) );
  OR2X1_RVT U6054 ( .A1(n12440), .A2(n5862), .Y(n6109) );
  OR2X1_RVT U6055 ( .A1(n5649), .A2(n5723), .Y(n6108) );
  OR2X1_RVT U6056 ( .A1(n316), .A2(n5680), .Y(n5723) );
  OR2X1_RVT U6057 ( .A1(n12443), .A2(n5841), .Y(n6104) );
  OR2X1_RVT U6058 ( .A1(n5716), .A2(n6110), .Y(n5841) );
  AND2X1_RVT U6059 ( .A1(n6111), .A2(n6112), .Y(n6103) );
  OR2X1_RVT U6060 ( .A1(n12412), .A2(n6113), .Y(n6112) );
  OR2X1_RVT U6061 ( .A1(n5719), .A2(n5668), .Y(n6111) );
  OR2X1_RVT U6062 ( .A1(n5642), .A2(n5927), .Y(n5668) );
  AND4X1_RVT U6063 ( .A1(n6115), .A2(n6116), .A3(n6117), .A4(n6118), .Y(n6114)
         );
  AND4X1_RVT U6064 ( .A1(n6119), .A2(n6120), .A3(n6121), .A4(n6122), .Y(n6118)
         );
  AND4X1_RVT U6065 ( .A1(n6123), .A2(n6124), .A3(n6125), .A4(n6126), .Y(n6122)
         );
  OR2X1_RVT U6066 ( .A1(n1391), .A2(n6127), .Y(n6121) );
  OR2X1_RVT U6067 ( .A1(n12203), .A2(n12194), .Y(n6127) );
  OR2X1_RVT U6068 ( .A1(n6128), .A2(n6129), .Y(n6120) );
  OR2X1_RVT U6069 ( .A1(n1325), .A2(n1388), .Y(n6129) );
  OR2X1_RVT U6070 ( .A1(n69), .A2(n6130), .Y(n6119) );
  OR2X1_RVT U6071 ( .A1(n6131), .A2(n6132), .Y(n6130) );
  AND4X1_RVT U6072 ( .A1(n6133), .A2(n6134), .A3(n6135), .A4(n6136), .Y(n6117)
         );
  OR2X1_RVT U6073 ( .A1(n6137), .A2(n12875), .Y(n6136) );
  AND2X1_RVT U6074 ( .A1(n6138), .A2(n6139), .Y(n6137) );
  AND2X1_RVT U6075 ( .A1(n6140), .A2(n6141), .Y(n6135) );
  OR2X1_RVT U6076 ( .A1(n6142), .A2(n6143), .Y(n6141) );
  AND2X1_RVT U6077 ( .A1(n1390), .A2(n1386), .Y(n6142) );
  OR2X1_RVT U6078 ( .A1(n6144), .A2(n12208), .Y(n6140) );
  AND2X1_RVT U6079 ( .A1(n1366), .A2(n6146), .Y(n6144) );
  OR2X1_RVT U6080 ( .A1(n6147), .A2(n1332), .Y(n6134) );
  AND2X1_RVT U6081 ( .A1(n6148), .A2(n6149), .Y(n6147) );
  AND2X1_RVT U6082 ( .A1(n6150), .A2(n6151), .Y(n6148) );
  AND2X1_RVT U6083 ( .A1(n6152), .A2(n6153), .Y(n6133) );
  OR2X1_RVT U6084 ( .A1(n6154), .A2(n12869), .Y(n6153) );
  AND2X1_RVT U6085 ( .A1(n6155), .A2(n6156), .Y(n6154) );
  OR2X1_RVT U6086 ( .A1(n6157), .A2(n12873), .Y(n6152) );
  AND2X1_RVT U6087 ( .A1(n6158), .A2(n6159), .Y(n6157) );
  AND4X1_RVT U6088 ( .A1(n6160), .A2(n6161), .A3(n6162), .A4(n6163), .Y(n6116)
         );
  AND4X1_RVT U6089 ( .A1(n6164), .A2(n6165), .A3(n6166), .A4(n6167), .Y(n6163)
         );
  OR2X1_RVT U6090 ( .A1(n6168), .A2(n12871), .Y(n6167) );
  AND2X1_RVT U6091 ( .A1(n6169), .A2(n6170), .Y(n6168) );
  OR2X1_RVT U6092 ( .A1(n6171), .A2(n12869), .Y(n6170) );
  AND2X1_RVT U6093 ( .A1(n6172), .A2(n6173), .Y(n6171) );
  OR2X1_RVT U6094 ( .A1(n1312), .A2(n12208), .Y(n6173) );
  AND2X1_RVT U6095 ( .A1(n6174), .A2(n6175), .Y(n6169) );
  OR2X1_RVT U6096 ( .A1(n12194), .A2(n6176), .Y(n6174) );
  OR2X1_RVT U6097 ( .A1(n6177), .A2(n12149), .Y(n6166) );
  AND2X1_RVT U6098 ( .A1(n6178), .A2(n6179), .Y(n6177) );
  OR2X1_RVT U6099 ( .A1(n1325), .A2(n6180), .Y(n6179) );
  AND2X1_RVT U6100 ( .A1(n6181), .A2(n6182), .Y(n6178) );
  OR2X1_RVT U6101 ( .A1(n12192), .A2(n6184), .Y(n6181) );
  OR2X1_RVT U6102 ( .A1(n6185), .A2(n1341), .Y(n6165) );
  AND4X1_RVT U6103 ( .A1(n6186), .A2(n6187), .A3(n6188), .A4(n6189), .Y(n6185)
         );
  OR2X1_RVT U6104 ( .A1(n1314), .A2(n6190), .Y(n6189) );
  AND2X1_RVT U6105 ( .A1(n6151), .A2(n6191), .Y(n6188) );
  OR2X1_RVT U6106 ( .A1(n12196), .A2(n6192), .Y(n6151) );
  OR2X1_RVT U6107 ( .A1(n6193), .A2(n12874), .Y(n6187) );
  AND2X1_RVT U6108 ( .A1(n6194), .A2(n6195), .Y(n6193) );
  OR2X1_RVT U6109 ( .A1(n12201), .A2(n12926), .Y(n6195) );
  OR2X1_RVT U6110 ( .A1(n12212), .A2(n12196), .Y(n6194) );
  OR2X1_RVT U6111 ( .A1(n12185), .A2(n6196), .Y(n6186) );
  OR2X1_RVT U6112 ( .A1(n6139), .A2(n1365), .Y(n6164) );
  OR2X1_RVT U6113 ( .A1(n6197), .A2(n76), .Y(n6162) );
  OR2X1_RVT U6114 ( .A1(n6198), .A2(n6199), .Y(n6161) );
  OR2X1_RVT U6115 ( .A1(n85), .A2(n6200), .Y(n6160) );
  AND4X1_RVT U6116 ( .A1(n6201), .A2(n6202), .A3(n6203), .A4(n6204), .Y(n6115)
         );
  OR2X1_RVT U6117 ( .A1(n12212), .A2(n6205), .Y(n6204) );
  AND2X1_RVT U6118 ( .A1(n6206), .A2(n6207), .Y(n6203) );
  OR2X1_RVT U6119 ( .A1(n12184), .A2(n6208), .Y(n6207) );
  OR2X1_RVT U6120 ( .A1(n12188), .A2(n6209), .Y(n6202) );
  AND2X1_RVT U6121 ( .A1(n6210), .A2(n6211), .Y(n6201) );
  OR2X1_RVT U6122 ( .A1(n12191), .A2(n1318), .Y(n6211) );
  OR2X1_RVT U6123 ( .A1(n1314), .A2(n6212), .Y(n1318) );
  OR2X1_RVT U6124 ( .A1(n73), .A2(n1325), .Y(n6212) );
  OR2X1_RVT U6125 ( .A1(n1307), .A2(n6213), .Y(n6210) );
  AND4X1_RVT U6126 ( .A1(n6215), .A2(n6216), .A3(n6217), .A4(n6218), .Y(n6214)
         );
  AND4X1_RVT U6127 ( .A1(n6219), .A2(n6220), .A3(n6221), .A4(n6222), .Y(n6218)
         );
  AND4X1_RVT U6128 ( .A1(n5855), .A2(n6045), .A3(n6223), .A4(n6224), .Y(n6222)
         );
  OR2X1_RVT U6129 ( .A1(n6225), .A2(n6226), .Y(n6045) );
  OR2X1_RVT U6130 ( .A1(n5640), .A2(n5910), .Y(n5855) );
  OR2X1_RVT U6131 ( .A1(n12686), .A2(n12428), .Y(n5910) );
  AND4X1_RVT U6132 ( .A1(n6113), .A2(n5979), .A3(n6102), .A4(n5637), .Y(n6221)
         );
  OR2X1_RVT U6133 ( .A1(n6227), .A2(n5827), .Y(n5637) );
  OR2X1_RVT U6134 ( .A1(n5642), .A2(n6228), .Y(n6102) );
  OR2X1_RVT U6135 ( .A1(n5675), .A2(n314), .Y(n5979) );
  OR2X1_RVT U6136 ( .A1(n5666), .A2(n6229), .Y(n6113) );
  OR2X1_RVT U6137 ( .A1(n12418), .A2(n12438), .Y(n6229) );
  AND4X1_RVT U6138 ( .A1(n6230), .A2(n6231), .A3(n6232), .A4(n6233), .Y(n6220)
         );
  OR2X1_RVT U6139 ( .A1(n5919), .A2(n6234), .Y(n6233) );
  OR2X1_RVT U6140 ( .A1(n12438), .A2(n5699), .Y(n6234) );
  OR2X1_RVT U6141 ( .A1(n5828), .A2(n6235), .Y(n6232) );
  OR2X1_RVT U6142 ( .A1(n12687), .A2(n5716), .Y(n6235) );
  OR2X1_RVT U6143 ( .A1(n6054), .A2(n6236), .Y(n6231) );
  OR2X1_RVT U6144 ( .A1(n6237), .A2(n5713), .Y(n6236) );
  OR2X1_RVT U6145 ( .A1(n12435), .A2(n6238), .Y(n6230) );
  OR2X1_RVT U6146 ( .A1(n6239), .A2(n12418), .Y(n6238) );
  AND2X1_RVT U6147 ( .A1(n5927), .A2(n6240), .Y(n6239) );
  AND2X1_RVT U6148 ( .A1(n6241), .A2(n6242), .Y(n6219) );
  OR2X1_RVT U6149 ( .A1(n6243), .A2(n5694), .Y(n6242) );
  AND2X1_RVT U6150 ( .A1(n6244), .A2(n6245), .Y(n6243) );
  OR2X1_RVT U6151 ( .A1(n12417), .A2(n5887), .Y(n6245) );
  OR2X1_RVT U6152 ( .A1(n12421), .A2(n5962), .Y(n6244) );
  AND2X1_RVT U6153 ( .A1(n6246), .A2(n6247), .Y(n6241) );
  OR2X1_RVT U6154 ( .A1(n6248), .A2(n5733), .Y(n6247) );
  AND2X1_RVT U6155 ( .A1(n6249), .A2(n6250), .Y(n6248) );
  OR2X1_RVT U6156 ( .A1(n12424), .A2(n324), .Y(n6250) );
  NAND2X1_RVT U6157 ( .A1(n5716), .A2(n12679), .Y(n6249) );
  OR2X1_RVT U6158 ( .A1(n6251), .A2(n316), .Y(n6246) );
  AND2X1_RVT U6159 ( .A1(n5940), .A2(n5817), .Y(n6251) );
  OR2X1_RVT U6160 ( .A1(n5666), .A2(n6252), .Y(n5817) );
  OR2X1_RVT U6161 ( .A1(n12690), .A2(n12413), .Y(n6252) );
  AND4X1_RVT U6162 ( .A1(n5834), .A2(n6253), .A3(n6026), .A4(n6254), .Y(n6217)
         );
  AND4X1_RVT U6163 ( .A1(n6255), .A2(n6256), .A3(n6257), .A4(n6258), .Y(n6254)
         );
  OR2X1_RVT U6164 ( .A1(n5797), .A2(n5718), .Y(n6258) );
  OR2X1_RVT U6165 ( .A1(n5735), .A2(n5764), .Y(n6257) );
  OR2X1_RVT U6166 ( .A1(n12678), .A2(n5989), .Y(n6256) );
  OR2X1_RVT U6167 ( .A1(n5713), .A2(n5695), .Y(n5989) );
  OR2X1_RVT U6168 ( .A1(n12686), .A2(n5777), .Y(n5695) );
  OR2X1_RVT U6169 ( .A1(n12427), .A2(n5818), .Y(n6255) );
  OR2X1_RVT U6170 ( .A1(n5699), .A2(n5927), .Y(n5818) );
  OR2X1_RVT U6171 ( .A1(n12411), .A2(n5903), .Y(n5927) );
  AND2X1_RVT U6172 ( .A1(n6259), .A2(n6260), .Y(n6026) );
  OR2X1_RVT U6173 ( .A1(n6261), .A2(n5766), .Y(n6260) );
  OR2X1_RVT U6174 ( .A1(n12437), .A2(n316), .Y(n6261) );
  OR2X1_RVT U6175 ( .A1(n6262), .A2(n5649), .Y(n6259) );
  OR2X1_RVT U6176 ( .A1(n12677), .A2(n5766), .Y(n5649) );
  OR2X1_RVT U6177 ( .A1(n5663), .A2(n5713), .Y(n6262) );
  OR2X1_RVT U6178 ( .A1(n12419), .A2(n6032), .Y(n6253) );
  AND2X1_RVT U6179 ( .A1(n6263), .A2(n6264), .Y(n5834) );
  OR2X1_RVT U6180 ( .A1(n5717), .A2(n5755), .Y(n6264) );
  OR2X1_RVT U6181 ( .A1(n6265), .A2(n6266), .Y(n6263) );
  AND4X1_RVT U6182 ( .A1(n6267), .A2(n6268), .A3(n6269), .A4(n6270), .Y(n6216)
         );
  OR2X1_RVT U6183 ( .A1(n6271), .A2(n5903), .Y(n6270) );
  AND2X1_RVT U6184 ( .A1(n6272), .A2(n5912), .Y(n6271) );
  OR2X1_RVT U6185 ( .A1(n12425), .A2(n6228), .Y(n5912) );
  OR2X1_RVT U6186 ( .A1(n6273), .A2(n12683), .Y(n6269) );
  AND2X1_RVT U6187 ( .A1(n5840), .A2(n5805), .Y(n6273) );
  OR2X1_RVT U6188 ( .A1(n12677), .A2(n5781), .Y(n5805) );
  OR2X1_RVT U6189 ( .A1(n6274), .A2(n5860), .Y(n6268) );
  AND2X1_RVT U6190 ( .A1(n6275), .A2(n6276), .Y(n6274) );
  OR2X1_RVT U6191 ( .A1(n12414), .A2(n5719), .Y(n6276) );
  AND2X1_RVT U6192 ( .A1(n6277), .A2(n5757), .Y(n6275) );
  OR2X1_RVT U6193 ( .A1(n314), .A2(n5716), .Y(n6277) );
  OR2X1_RVT U6194 ( .A1(n6278), .A2(n5657), .Y(n6267) );
  AND2X1_RVT U6195 ( .A1(n6279), .A2(n6280), .Y(n6278) );
  NAND2X1_RVT U6196 ( .A1(n5642), .A2(n6020), .Y(n6280) );
  AND2X1_RVT U6197 ( .A1(n6281), .A2(n5870), .Y(n6279) );
  OR2X1_RVT U6198 ( .A1(n5803), .A2(n6228), .Y(n5870) );
  OR2X1_RVT U6199 ( .A1(n12434), .A2(n6282), .Y(n6281) );
  AND4X1_RVT U6200 ( .A1(n6283), .A2(n6284), .A3(n6285), .A4(n6286), .Y(n6215)
         );
  OR2X1_RVT U6201 ( .A1(n6287), .A2(n5680), .Y(n6286) );
  AND2X1_RVT U6202 ( .A1(n6288), .A2(n5821), .Y(n6287) );
  AND2X1_RVT U6203 ( .A1(n6289), .A2(n5843), .Y(n6288) );
  OR2X1_RVT U6204 ( .A1(n316), .A2(n6266), .Y(n5843) );
  OR2X1_RVT U6205 ( .A1(n12413), .A2(n5777), .Y(n6266) );
  OR2X1_RVT U6206 ( .A1(n6290), .A2(n12430), .Y(n6285) );
  AND2X1_RVT U6207 ( .A1(n6291), .A2(n6292), .Y(n6290) );
  OR2X1_RVT U6208 ( .A1(n6293), .A2(n12675), .Y(n6292) );
  AND2X1_RVT U6209 ( .A1(n6294), .A2(n6295), .Y(n6293) );
  OR2X1_RVT U6210 ( .A1(n12412), .A2(n6054), .Y(n6295) );
  OR2X1_RVT U6211 ( .A1(n12682), .A2(n5700), .Y(n6294) );
  AND2X1_RVT U6212 ( .A1(n6296), .A2(n6297), .Y(n6291) );
  OR2X1_RVT U6213 ( .A1(n5666), .A2(n6298), .Y(n6296) );
  OR2X1_RVT U6214 ( .A1(n6299), .A2(n5700), .Y(n6284) );
  AND4X1_RVT U6215 ( .A1(n6300), .A2(n6301), .A3(n6302), .A4(n5666), .Y(n6299)
         );
  OR2X1_RVT U6216 ( .A1(n12683), .A2(n5716), .Y(n6302) );
  OR2X1_RVT U6217 ( .A1(n12424), .A2(n5735), .Y(n6301) );
  OR2X1_RVT U6218 ( .A1(n5788), .A2(n5766), .Y(n6300) );
  OR2X1_RVT U6219 ( .A1(n6303), .A2(n5642), .Y(n6283) );
  AND4X1_RVT U6220 ( .A1(n6067), .A2(n6304), .A3(n5865), .A4(n5781), .Y(n6303)
         );
  OR2X1_RVT U6221 ( .A1(n5735), .A2(n6298), .Y(n5865) );
  OR2X1_RVT U6222 ( .A1(n5903), .A2(n6110), .Y(n6304) );
  OR2X1_RVT U6223 ( .A1(n12418), .A2(n5868), .Y(n6067) );
  AND4X1_RVT U6224 ( .A1(n6306), .A2(n6307), .A3(n6308), .A4(n6309), .Y(n6305)
         );
  AND4X1_RVT U6225 ( .A1(n5718), .A2(n5954), .A3(n6310), .A4(n6311), .Y(n6309)
         );
  AND4X1_RVT U6226 ( .A1(n6033), .A2(n5978), .A3(n6223), .A4(n6224), .Y(n6311)
         );
  OR2X1_RVT U6227 ( .A1(n6226), .A2(n5639), .Y(n6224) );
  OR2X1_RVT U6228 ( .A1(n12681), .A2(n5757), .Y(n5639) );
  OR2X1_RVT U6229 ( .A1(n5656), .A2(n6265), .Y(n6223) );
  OR2X1_RVT U6230 ( .A1(n12686), .A2(n12432), .Y(n6265) );
  OR2X1_RVT U6231 ( .A1(n12675), .A2(n5777), .Y(n5656) );
  OR2X1_RVT U6232 ( .A1(n12687), .A2(n5675), .Y(n5978) );
  OR2X1_RVT U6233 ( .A1(n12441), .A2(n12425), .Y(n5675) );
  OR2X1_RVT U6234 ( .A1(n5797), .A2(n6312), .Y(n6033) );
  OR2X1_RVT U6235 ( .A1(n12432), .A2(n5701), .Y(n6312) );
  OR2X1_RVT U6236 ( .A1(n5699), .A2(n6313), .Y(n6310) );
  OR2X1_RVT U6237 ( .A1(n5827), .A2(n12423), .Y(n6313) );
  OR2X1_RVT U6238 ( .A1(n5766), .A2(n6314), .Y(n5954) );
  OR2X1_RVT U6239 ( .A1(n5700), .A2(n12430), .Y(n6314) );
  OR2X1_RVT U6240 ( .A1(n12679), .A2(n6225), .Y(n5718) );
  OR2X1_RVT U6241 ( .A1(n12425), .A2(n5717), .Y(n6225) );
  AND4X1_RVT U6242 ( .A1(n6315), .A2(n6316), .A3(n6317), .A4(n6318), .Y(n6308)
         );
  AND4X1_RVT U6243 ( .A1(n6319), .A2(n6320), .A3(n6321), .A4(n6322), .Y(n6318)
         );
  OR2X1_RVT U6244 ( .A1(n5733), .A2(n6323), .Y(n6322) );
  OR2X1_RVT U6245 ( .A1(n12414), .A2(n5803), .Y(n6323) );
  OR2X1_RVT U6246 ( .A1(n5716), .A2(n6324), .Y(n6321) );
  OR2X1_RVT U6247 ( .A1(n6325), .A2(n5680), .Y(n6324) );
  AND2X1_RVT U6248 ( .A1(n5659), .A2(n5719), .Y(n6325) );
  OR2X1_RVT U6249 ( .A1(n6326), .A2(n6327), .Y(n6320) );
  AND2X1_RVT U6250 ( .A1(n5874), .A2(n5830), .Y(n6326) );
  OR2X1_RVT U6251 ( .A1(n12680), .A2(n324), .Y(n5830) );
  OR2X1_RVT U6252 ( .A1(n12676), .A2(n12435), .Y(n5874) );
  OR2X1_RVT U6253 ( .A1(n6328), .A2(n5714), .Y(n6319) );
  AND2X1_RVT U6254 ( .A1(n6110), .A2(n6329), .Y(n6328) );
  OR2X1_RVT U6255 ( .A1(n12678), .A2(n316), .Y(n6329) );
  OR2X1_RVT U6256 ( .A1(n6330), .A2(n12437), .Y(n6317) );
  AND2X1_RVT U6257 ( .A1(n6101), .A2(n6331), .Y(n6330) );
  OR2X1_RVT U6258 ( .A1(n5707), .A2(n6054), .Y(n6331) );
  OR2X1_RVT U6259 ( .A1(n12418), .A2(n5919), .Y(n6101) );
  OR2X1_RVT U6260 ( .A1(n12682), .A2(n5707), .Y(n5919) );
  OR2X1_RVT U6261 ( .A1(n6332), .A2(n5868), .Y(n6316) );
  AND2X1_RVT U6262 ( .A1(n5821), .A2(n6093), .Y(n6332) );
  OR2X1_RVT U6263 ( .A1(n5677), .A2(n5766), .Y(n5821) );
  OR2X1_RVT U6264 ( .A1(n6333), .A2(n5757), .Y(n6315) );
  AND2X1_RVT U6265 ( .A1(n5720), .A2(n5722), .Y(n6333) );
  AND4X1_RVT U6266 ( .A1(n6334), .A2(n6335), .A3(n6336), .A4(n6337), .Y(n6307)
         );
  AND4X1_RVT U6267 ( .A1(n6338), .A2(n6339), .A3(n6340), .A4(n6341), .Y(n6337)
         );
  OR2X1_RVT U6268 ( .A1(n6342), .A2(n12421), .Y(n6341) );
  AND2X1_RVT U6269 ( .A1(n5648), .A2(n5940), .Y(n6342) );
  OR2X1_RVT U6270 ( .A1(n5797), .A2(n5828), .Y(n5940) );
  OR2X1_RVT U6271 ( .A1(n12424), .A2(n5680), .Y(n5828) );
  OR2X1_RVT U6272 ( .A1(n12428), .A2(n6343), .Y(n5648) );
  OR2X1_RVT U6273 ( .A1(n12411), .A2(n12417), .Y(n6343) );
  OR2X1_RVT U6274 ( .A1(n6344), .A2(n12435), .Y(n6340) );
  AND2X1_RVT U6275 ( .A1(n5957), .A2(n6345), .Y(n6344) );
  OR2X1_RVT U6276 ( .A1(n12440), .A2(n314), .Y(n6345) );
  OR2X1_RVT U6277 ( .A1(n12438), .A2(n5764), .Y(n5957) );
  OR2X1_RVT U6278 ( .A1(n6346), .A2(n12416), .Y(n6339) );
  AND2X1_RVT U6279 ( .A1(n5975), .A2(n6347), .Y(n6346) );
  OR2X1_RVT U6280 ( .A1(n12441), .A2(n5700), .Y(n6347) );
  OR2X1_RVT U6281 ( .A1(n5642), .A2(n6348), .Y(n5975) );
  OR2X1_RVT U6282 ( .A1(n6349), .A2(n5701), .Y(n6338) );
  AND2X1_RVT U6283 ( .A1(n6350), .A2(n6351), .Y(n6349) );
  OR2X1_RVT U6284 ( .A1(n5757), .A2(n12438), .Y(n6351) );
  AND2X1_RVT U6285 ( .A1(n6352), .A2(n5733), .Y(n6350) );
  OR2X1_RVT U6286 ( .A1(n5719), .A2(n5680), .Y(n5733) );
  OR2X1_RVT U6287 ( .A1(n12413), .A2(n5764), .Y(n6352) );
  OR2X1_RVT U6288 ( .A1(n12690), .A2(n5719), .Y(n5764) );
  OR2X1_RVT U6289 ( .A1(n6353), .A2(n5777), .Y(n6336) );
  AND4X1_RVT U6290 ( .A1(n6354), .A2(n6355), .A3(n5930), .A4(n5840), .Y(n6353)
         );
  OR2X1_RVT U6291 ( .A1(n5903), .A2(n6003), .Y(n5840) );
  OR2X1_RVT U6292 ( .A1(n5735), .A2(n6282), .Y(n5930) );
  OR2X1_RVT U6293 ( .A1(n12419), .A2(n12412), .Y(n6282) );
  OR2X1_RVT U6294 ( .A1(n316), .A2(n5657), .Y(n6355) );
  OR2X1_RVT U6295 ( .A1(n314), .A2(n12438), .Y(n6354) );
  OR2X1_RVT U6296 ( .A1(n6356), .A2(n5713), .Y(n6335) );
  AND2X1_RVT U6297 ( .A1(n6357), .A2(n5734), .Y(n6356) );
  AND2X1_RVT U6298 ( .A1(n6289), .A2(n5984), .Y(n6357) );
  OR2X1_RVT U6299 ( .A1(n6358), .A2(n12687), .Y(n5984) );
  AND2X1_RVT U6300 ( .A1(n5755), .A2(n6359), .Y(n6358) );
  OR2X1_RVT U6301 ( .A1(n12416), .A2(n5642), .Y(n6359) );
  OR2X1_RVT U6302 ( .A1(n5803), .A2(n5941), .Y(n6289) );
  OR2X1_RVT U6303 ( .A1(n5788), .A2(n5677), .Y(n5941) );
  OR2X1_RVT U6304 ( .A1(n6360), .A2(n5781), .Y(n6334) );
  AND2X1_RVT U6305 ( .A1(n6361), .A2(n12424), .Y(n6360) );
  AND2X1_RVT U6306 ( .A1(n6362), .A2(n5962), .Y(n6361) );
  OR2X1_RVT U6307 ( .A1(n5803), .A2(n5903), .Y(n6362) );
  AND4X1_RVT U6308 ( .A1(n6363), .A2(n6364), .A3(n6365), .A4(n6366), .Y(n6306)
         );
  AND2X1_RVT U6309 ( .A1(n6367), .A2(n6368), .Y(n6366) );
  OR2X1_RVT U6310 ( .A1(n12683), .A2(n5883), .Y(n6368) );
  OR2X1_RVT U6311 ( .A1(n12432), .A2(n6369), .Y(n5883) );
  OR2X1_RVT U6312 ( .A1(n5699), .A2(n5788), .Y(n6369) );
  AND2X1_RVT U6313 ( .A1(n6370), .A2(n6371), .Y(n6367) );
  OR2X1_RVT U6314 ( .A1(n5672), .A2(n5683), .Y(n6371) );
  OR2X1_RVT U6315 ( .A1(n5716), .A2(n5911), .Y(n5683) );
  OR2X1_RVT U6316 ( .A1(n12679), .A2(n5677), .Y(n5911) );
  OR2X1_RVT U6317 ( .A1(n5719), .A2(n5796), .Y(n6370) );
  OR2X1_RVT U6318 ( .A1(n5707), .A2(n6372), .Y(n5796) );
  OR2X1_RVT U6319 ( .A1(n5707), .A2(n5887), .Y(n6365) );
  OR2X1_RVT U6320 ( .A1(n316), .A2(n12434), .Y(n5887) );
  OR2X1_RVT U6321 ( .A1(n6373), .A2(n5663), .Y(n6364) );
  AND4X1_RVT U6322 ( .A1(n6374), .A2(n6375), .A3(n6376), .A4(n6377), .Y(n6373)
         );
  OR2X1_RVT U6323 ( .A1(n12677), .A2(n6378), .Y(n6376) );
  OR2X1_RVT U6324 ( .A1(n6379), .A2(n12684), .Y(n6378) );
  AND2X1_RVT U6325 ( .A1(n5714), .A2(n6380), .Y(n6379) );
  OR2X1_RVT U6326 ( .A1(n12427), .A2(n6381), .Y(n6375) );
  OR2X1_RVT U6327 ( .A1(n6020), .A2(n5657), .Y(n6381) );
  OR2X1_RVT U6328 ( .A1(n5640), .A2(n5666), .Y(n6374) );
  OR2X1_RVT U6329 ( .A1(n12681), .A2(n5766), .Y(n5666) );
  OR2X1_RVT U6330 ( .A1(n6240), .A2(n6054), .Y(n6363) );
  OR2X1_RVT U6331 ( .A1(n12443), .A2(n5677), .Y(n6054) );
  AND4X1_RVT U6332 ( .A1(n6383), .A2(n6384), .A3(n6385), .A4(n6386), .Y(n6382)
         );
  AND4X1_RVT U6333 ( .A1(n6387), .A2(n6388), .A3(n6389), .A4(n6390), .Y(n6386)
         );
  AND4X1_RVT U6334 ( .A1(n6391), .A2(n6392), .A3(n6393), .A4(n6394), .Y(n6390)
         );
  OR2X1_RVT U6335 ( .A1(n6228), .A2(n6372), .Y(n6394) );
  OR2X1_RVT U6336 ( .A1(n12680), .A2(n12437), .Y(n6372) );
  OR2X1_RVT U6337 ( .A1(n12411), .A2(n12421), .Y(n6228) );
  OR2X1_RVT U6338 ( .A1(n6395), .A2(n5714), .Y(n6393) );
  AND2X1_RVT U6339 ( .A1(n5660), .A2(n6327), .Y(n6395) );
  OR2X1_RVT U6340 ( .A1(n316), .A2(n6396), .Y(n5660) );
  OR2X1_RVT U6341 ( .A1(n12411), .A2(n12677), .Y(n6396) );
  OR2X1_RVT U6342 ( .A1(n6397), .A2(n5642), .Y(n6392) );
  OR2X1_RVT U6343 ( .A1(n12425), .A2(n5803), .Y(n5642) );
  AND2X1_RVT U6344 ( .A1(n5778), .A2(n6398), .Y(n6397) );
  OR2X1_RVT U6345 ( .A1(n5657), .A2(n5859), .Y(n6398) );
  OR2X1_RVT U6346 ( .A1(n12429), .A2(n12417), .Y(n5657) );
  OR2X1_RVT U6347 ( .A1(n5903), .A2(n6399), .Y(n5778) );
  OR2X1_RVT U6348 ( .A1(n12688), .A2(n12432), .Y(n6399) );
  OR2X1_RVT U6349 ( .A1(n6400), .A2(n5701), .Y(n6391) );
  AND2X1_RVT U6350 ( .A1(n6098), .A2(n6401), .Y(n6400) );
  OR2X1_RVT U6351 ( .A1(n6402), .A2(n12677), .Y(n6401) );
  AND2X1_RVT U6352 ( .A1(n5757), .A2(n6110), .Y(n6402) );
  OR2X1_RVT U6353 ( .A1(n12685), .A2(n5719), .Y(n6110) );
  OR2X1_RVT U6354 ( .A1(n12438), .A2(n6403), .Y(n6098) );
  OR2X1_RVT U6355 ( .A1(n12690), .A2(n12686), .Y(n6403) );
  OR2X1_RVT U6356 ( .A1(n6404), .A2(n12416), .Y(n6389) );
  AND2X1_RVT U6357 ( .A1(n6405), .A2(n6406), .Y(n6404) );
  OR2X1_RVT U6358 ( .A1(n6407), .A2(n5803), .Y(n6406) );
  AND2X1_RVT U6359 ( .A1(n5868), .A2(n6408), .Y(n6407) );
  OR2X1_RVT U6360 ( .A1(n5659), .A2(n5781), .Y(n6405) );
  OR2X1_RVT U6361 ( .A1(n12430), .A2(n5717), .Y(n5781) );
  OR2X1_RVT U6362 ( .A1(n6409), .A2(n12686), .Y(n6388) );
  AND2X1_RVT U6363 ( .A1(n5873), .A2(n6032), .Y(n6409) );
  OR2X1_RVT U6364 ( .A1(n12428), .A2(n6410), .Y(n6032) );
  OR2X1_RVT U6365 ( .A1(n5713), .A2(n12417), .Y(n6410) );
  OR2X1_RVT U6366 ( .A1(n5659), .A2(n6240), .Y(n5873) );
  OR2X1_RVT U6367 ( .A1(n12417), .A2(n12432), .Y(n6240) );
  OR2X1_RVT U6368 ( .A1(n6411), .A2(n12414), .Y(n6387) );
  AND2X1_RVT U6369 ( .A1(n5913), .A2(n6412), .Y(n6411) );
  OR2X1_RVT U6370 ( .A1(n6227), .A2(n5707), .Y(n6412) );
  OR2X1_RVT U6371 ( .A1(n5766), .A2(n6348), .Y(n5913) );
  OR2X1_RVT U6372 ( .A1(n12685), .A2(n316), .Y(n6348) );
  AND2X1_RVT U6373 ( .A1(n12418), .A2(n12688), .Y(n6009) );
  AND4X1_RVT U6374 ( .A1(n6413), .A2(n6414), .A3(n6415), .A4(n6416), .Y(n6385)
         );
  AND4X1_RVT U6375 ( .A1(n6417), .A2(n6418), .A3(n6419), .A4(n6420), .Y(n6416)
         );
  OR2X1_RVT U6376 ( .A1(n6421), .A2(n12423), .Y(n6420) );
  AND2X1_RVT U6377 ( .A1(n5900), .A2(n5971), .Y(n6421) );
  OR2X1_RVT U6378 ( .A1(n5716), .A2(n6327), .Y(n5971) );
  OR2X1_RVT U6379 ( .A1(n12688), .A2(n5713), .Y(n6327) );
  OR2X1_RVT U6380 ( .A1(n12675), .A2(n12413), .Y(n5716) );
  OR2X1_RVT U6381 ( .A1(n12414), .A2(n6003), .Y(n5900) );
  OR2X1_RVT U6382 ( .A1(n12418), .A2(n12432), .Y(n6003) );
  OR2X1_RVT U6383 ( .A1(n6422), .A2(n12684), .Y(n6419) );
  AND2X1_RVT U6384 ( .A1(n6062), .A2(n6423), .Y(n6422) );
  OR2X1_RVT U6385 ( .A1(n6020), .A2(n5730), .Y(n6423) );
  OR2X1_RVT U6386 ( .A1(n5903), .A2(n6424), .Y(n5730) );
  OR2X1_RVT U6387 ( .A1(n12443), .A2(n12419), .Y(n6424) );
  OR2X1_RVT U6388 ( .A1(n12427), .A2(n6425), .Y(n6062) );
  OR2X1_RVT U6389 ( .A1(n5903), .A2(n5699), .Y(n6425) );
  OR2X1_RVT U6390 ( .A1(n6426), .A2(n12690), .Y(n6418) );
  AND2X1_RVT U6391 ( .A1(n6008), .A2(n5937), .Y(n6426) );
  OR2X1_RVT U6392 ( .A1(n5719), .A2(n5755), .Y(n5937) );
  OR2X1_RVT U6393 ( .A1(n12682), .A2(n5903), .Y(n5755) );
  OR2X1_RVT U6394 ( .A1(n6227), .A2(n5735), .Y(n6008) );
  OR2X1_RVT U6395 ( .A1(n12424), .A2(n12687), .Y(n6227) );
  OR2X1_RVT U6396 ( .A1(n6427), .A2(n5777), .Y(n6417) );
  AND2X1_RVT U6397 ( .A1(n6428), .A2(n6429), .Y(n6427) );
  OR2X1_RVT U6398 ( .A1(n5699), .A2(n6226), .Y(n6429) );
  OR2X1_RVT U6399 ( .A1(n12684), .A2(n324), .Y(n6226) );
  AND2X1_RVT U6400 ( .A1(n6430), .A2(n5994), .Y(n6428) );
  OR2X1_RVT U6401 ( .A1(n5707), .A2(n6431), .Y(n5994) );
  OR2X1_RVT U6402 ( .A1(n12440), .A2(n12419), .Y(n6431) );
  OR2X1_RVT U6403 ( .A1(n5763), .A2(n5700), .Y(n6415) );
  OR2X1_RVT U6404 ( .A1(n12677), .A2(n5659), .Y(n5763) );
  OR2X1_RVT U6405 ( .A1(n6432), .A2(n5663), .Y(n6414) );
  AND2X1_RVT U6406 ( .A1(n6433), .A2(n5844), .Y(n6432) );
  AND2X1_RVT U6407 ( .A1(n6434), .A2(n6435), .Y(n5844) );
  OR2X1_RVT U6408 ( .A1(n12428), .A2(n5868), .Y(n6435) );
  OR2X1_RVT U6409 ( .A1(n5766), .A2(n5640), .Y(n6434) );
  OR2X1_RVT U6410 ( .A1(n12413), .A2(n5713), .Y(n5640) );
  AND2X1_RVT U6411 ( .A1(n6436), .A2(n6030), .Y(n6433) );
  OR2X1_RVT U6412 ( .A1(n5797), .A2(n6380), .Y(n6030) );
  OR2X1_RVT U6413 ( .A1(n12679), .A2(n314), .Y(n6380) );
  OR2X1_RVT U6414 ( .A1(n5659), .A2(n5826), .Y(n6436) );
  OR2X1_RVT U6415 ( .A1(n12412), .A2(n6437), .Y(n5826) );
  OR2X1_RVT U6416 ( .A1(n12675), .A2(n12441), .Y(n6437) );
  OR2X1_RVT U6417 ( .A1(n6438), .A2(n12675), .Y(n6413) );
  AND4X1_RVT U6418 ( .A1(n6439), .A2(n6440), .A3(n6441), .A4(n6272), .Y(n6438)
         );
  OR2X1_RVT U6419 ( .A1(n5713), .A2(n6093), .Y(n6272) );
  OR2X1_RVT U6420 ( .A1(n12680), .A2(n12686), .Y(n6093) );
  OR2X1_RVT U6421 ( .A1(n5713), .A2(n6442), .Y(n6441) );
  OR2X1_RVT U6422 ( .A1(n12418), .A2(n12423), .Y(n6442) );
  OR2X1_RVT U6423 ( .A1(n12685), .A2(n5672), .Y(n5713) );
  OR2X1_RVT U6424 ( .A1(n6443), .A2(n5794), .Y(n6440) );
  OR2X1_RVT U6425 ( .A1(n12412), .A2(n5638), .Y(n5794) );
  AND2X1_RVT U6426 ( .A1(n5777), .A2(n6444), .Y(n6443) );
  OR2X1_RVT U6427 ( .A1(n12683), .A2(n5677), .Y(n6444) );
  OR2X1_RVT U6428 ( .A1(n12679), .A2(n12423), .Y(n5777) );
  OR2X1_RVT U6429 ( .A1(n12681), .A2(n6408), .Y(n6439) );
  OR2X1_RVT U6430 ( .A1(n12685), .A2(n5717), .Y(n6408) );
  OR2X1_RVT U6431 ( .A1(n5663), .A2(n314), .Y(n5717) );
  AND4X1_RVT U6432 ( .A1(n6445), .A2(n6446), .A3(n6447), .A4(n6448), .Y(n6384)
         );
  AND4X1_RVT U6433 ( .A1(n6449), .A2(n6450), .A3(n6451), .A4(n6452), .Y(n6448)
         );
  OR2X1_RVT U6434 ( .A1(n5735), .A2(n5862), .Y(n6452) );
  OR2X1_RVT U6435 ( .A1(n12425), .A2(n5757), .Y(n5862) );
  OR2X1_RVT U6436 ( .A1(n12429), .A2(n5903), .Y(n5735) );
  OR2X1_RVT U6437 ( .A1(n5722), .A2(n6298), .Y(n6451) );
  OR2X1_RVT U6438 ( .A1(n12689), .A2(n12412), .Y(n6298) );
  OR2X1_RVT U6439 ( .A1(n5788), .A2(n5714), .Y(n5722) );
  OR2X1_RVT U6440 ( .A1(n5707), .A2(n5734), .Y(n6450) );
  OR2X1_RVT U6441 ( .A1(n12421), .A2(n12434), .Y(n5734) );
  OR2X1_RVT U6442 ( .A1(n12411), .A2(n12676), .Y(n5707) );
  OR2X1_RVT U6443 ( .A1(n324), .A2(n6073), .Y(n6449) );
  OR2X1_RVT U6444 ( .A1(n12419), .A2(n5860), .Y(n6073) );
  OR2X1_RVT U6445 ( .A1(n5677), .A2(n6107), .Y(n6447) );
  OR2X1_RVT U6446 ( .A1(n324), .A2(n6453), .Y(n6107) );
  OR2X1_RVT U6447 ( .A1(n12682), .A2(n12432), .Y(n6453) );
  AND2X1_RVT U6448 ( .A1(n12413), .A2(n12416), .Y(n6237) );
  OR2X1_RVT U6449 ( .A1(n5719), .A2(n5667), .Y(n6446) );
  OR2X1_RVT U6450 ( .A1(n12441), .A2(n6454), .Y(n5667) );
  OR2X1_RVT U6451 ( .A1(n12683), .A2(n12675), .Y(n6454) );
  OR2X1_RVT U6452 ( .A1(n12418), .A2(n5699), .Y(n5719) );
  OR2X1_RVT U6453 ( .A1(n5766), .A2(n6430), .Y(n6445) );
  OR2X1_RVT U6454 ( .A1(n12414), .A2(n5721), .Y(n6430) );
  OR2X1_RVT U6455 ( .A1(n12685), .A2(n12686), .Y(n5721) );
  AND4X1_RVT U6456 ( .A1(n6455), .A2(n5832), .A3(n6456), .A4(n6457), .Y(n6383)
         );
  OR2X1_RVT U6457 ( .A1(n12418), .A2(n6377), .Y(n6457) );
  OR2X1_RVT U6458 ( .A1(n12681), .A2(n5827), .Y(n6377) );
  OR2X1_RVT U6459 ( .A1(n12416), .A2(n5868), .Y(n5827) );
  OR2X1_RVT U6460 ( .A1(n12411), .A2(n5694), .Y(n5868) );
  AND2X1_RVT U6461 ( .A1(n6458), .A2(n6459), .Y(n6456) );
  OR2X1_RVT U6462 ( .A1(n12440), .A2(n6297), .Y(n6459) );
  OR2X1_RVT U6463 ( .A1(n5766), .A2(n5859), .Y(n6297) );
  OR2X1_RVT U6464 ( .A1(n12418), .A2(n12412), .Y(n5859) );
  OR2X1_RVT U6465 ( .A1(n12413), .A2(n5655), .Y(n5694) );
  OR2X1_RVT U6466 ( .A1(n12688), .A2(n5928), .Y(n6458) );
  OR2X1_RVT U6467 ( .A1(n12437), .A2(n5962), .Y(n5928) );
  OR2X1_RVT U6468 ( .A1(n12680), .A2(n12675), .Y(n5962) );
  OR2X1_RVT U6469 ( .A1(n12678), .A2(n12429), .Y(n5638) );
  AND2X1_RVT U6470 ( .A1(n6460), .A2(n6461), .Y(n5832) );
  OR2X1_RVT U6471 ( .A1(n5714), .A2(n5700), .Y(n6461) );
  OR2X1_RVT U6472 ( .A1(n12687), .A2(n5672), .Y(n5700) );
  AND2X1_RVT U6473 ( .A1(n5699), .A2(n5663), .Y(n5752) );
  OR2X1_RVT U6474 ( .A1(n12424), .A2(n5766), .Y(n5714) );
  OR2X1_RVT U6475 ( .A1(n12676), .A2(n5803), .Y(n5766) );
  OR2X1_RVT U6476 ( .A1(n6462), .A2(n5757), .Y(n6460) );
  OR2X1_RVT U6477 ( .A1(n12418), .A2(n314), .Y(n5757) );
  AND2X1_RVT U6478 ( .A1(n12689), .A2(n12411), .Y(n6020) );
  OR2X1_RVT U6479 ( .A1(n12417), .A2(n5860), .Y(n6462) );
  OR2X1_RVT U6480 ( .A1(n12685), .A2(n12434), .Y(n5860) );
  AND2X1_RVT U6481 ( .A1(n6463), .A2(n6464), .Y(n6455) );
  OR2X1_RVT U6482 ( .A1(n5680), .A2(n6013), .Y(n6464) );
  OR2X1_RVT U6483 ( .A1(n12419), .A2(n5720), .Y(n6013) );
  OR2X1_RVT U6484 ( .A1(n12434), .A2(n5797), .Y(n5720) );
  OR2X1_RVT U6485 ( .A1(n12414), .A2(n12417), .Y(n5797) );
  OR2X1_RVT U6486 ( .A1(n12682), .A2(n12680), .Y(n5659) );
  OR2X1_RVT U6487 ( .A1(n12690), .A2(n12684), .Y(n5680) );
  XOR2X1_RVT U6488 ( .A1(key[4]), .A2(state[4]), .Y(n5655) );
  OR2X1_RVT U6489 ( .A1(n5672), .A2(n5801), .Y(n6463) );
  OR2X1_RVT U6490 ( .A1(n5903), .A2(n6094), .Y(n5801) );
  OR2X1_RVT U6491 ( .A1(n12421), .A2(n5701), .Y(n6094) );
  OR2X1_RVT U6492 ( .A1(n12683), .A2(n5803), .Y(n5701) );
  XOR2X1_RVT U6493 ( .A1(key[2]), .A2(state[2]), .Y(n5803) );
  XOR2X1_RVT U6494 ( .A1(key[3]), .A2(state[3]), .Y(n5737) );
  OR2X1_RVT U6495 ( .A1(n12688), .A2(n12419), .Y(n5677) );
  XOR2X1_RVT U6496 ( .A1(key[5]), .A2(state[5]), .Y(n5663) );
  XOR2X1_RVT U6497 ( .A1(key[6]), .A2(state[6]), .Y(n5699) );
  OR2X1_RVT U6498 ( .A1(n12678), .A2(n12417), .Y(n5903) );
  XOR2X1_RVT U6499 ( .A1(key[0]), .A2(state[0]), .Y(n5678) );
  XOR2X1_RVT U6500 ( .A1(key[1]), .A2(state[1]), .Y(n5788) );
  XOR2X1_RVT U6501 ( .A1(key[7]), .A2(state[7]), .Y(n5672) );
  AND4X1_RVT U6502 ( .A1(n6466), .A2(n6467), .A3(n6468), .A4(n6469), .Y(n6465)
         );
  AND4X1_RVT U6503 ( .A1(n6470), .A2(n6471), .A3(n6472), .A4(n6473), .Y(n6469)
         );
  AND4X1_RVT U6504 ( .A1(n6474), .A2(n6475), .A3(n6476), .A4(n6477), .Y(n6473)
         );
  OR2X1_RVT U6505 ( .A1(n12405), .A2(n6479), .Y(n6472) );
  OR2X1_RVT U6506 ( .A1(n6480), .A2(n6481), .Y(n6470) );
  OR2X1_RVT U6507 ( .A1(n12800), .A2(n6482), .Y(n6481) );
  AND4X1_RVT U6508 ( .A1(n6483), .A2(n6484), .A3(n6485), .A4(n6486), .Y(n6468)
         );
  OR2X1_RVT U6509 ( .A1(n6487), .A2(n12798), .Y(n6486) );
  AND2X1_RVT U6510 ( .A1(n6488), .A2(n6489), .Y(n6487) );
  AND2X1_RVT U6511 ( .A1(n6490), .A2(n6491), .Y(n6485) );
  OR2X1_RVT U6512 ( .A1(n6492), .A2(n176), .Y(n6491) );
  AND2X1_RVT U6513 ( .A1(n6493), .A2(n6494), .Y(n6492) );
  OR2X1_RVT U6514 ( .A1(n12396), .A2(n6496), .Y(n6494) );
  OR2X1_RVT U6515 ( .A1(n6482), .A2(n6497), .Y(n6493) );
  OR2X1_RVT U6516 ( .A1(n6498), .A2(n12402), .Y(n6490) );
  AND2X1_RVT U6517 ( .A1(n6500), .A2(n6501), .Y(n6498) );
  OR2X1_RVT U6518 ( .A1(n6502), .A2(n6503), .Y(n6484) );
  AND2X1_RVT U6519 ( .A1(n6504), .A2(n6505), .Y(n6502) );
  OR2X1_RVT U6520 ( .A1(n12397), .A2(n6506), .Y(n6505) );
  AND2X1_RVT U6521 ( .A1(n6507), .A2(n6508), .Y(n6504) );
  AND2X1_RVT U6522 ( .A1(n6509), .A2(n6510), .Y(n6483) );
  OR2X1_RVT U6523 ( .A1(n6511), .A2(n12379), .Y(n6510) );
  AND2X1_RVT U6524 ( .A1(n6513), .A2(n6514), .Y(n6511) );
  OR2X1_RVT U6525 ( .A1(n6515), .A2(n6516), .Y(n6514) );
  OR2X1_RVT U6526 ( .A1(n12388), .A2(n12383), .Y(n6516) );
  OR2X1_RVT U6527 ( .A1(n6519), .A2(n6520), .Y(n6509) );
  AND2X1_RVT U6528 ( .A1(n6521), .A2(n6522), .Y(n6519) );
  AND2X1_RVT U6529 ( .A1(n6523), .A2(n6524), .Y(n6521) );
  AND4X1_RVT U6530 ( .A1(n6525), .A2(n6526), .A3(n6527), .A4(n6528), .Y(n6467)
         );
  AND4X1_RVT U6531 ( .A1(n6529), .A2(n6530), .A3(n6531), .A4(n6532), .Y(n6528)
         );
  OR2X1_RVT U6532 ( .A1(n6533), .A2(n12408), .Y(n6532) );
  AND4X1_RVT U6533 ( .A1(n6535), .A2(n6536), .A3(n6537), .A4(n6538), .Y(n6533)
         );
  OR2X1_RVT U6534 ( .A1(n6539), .A2(n6506), .Y(n6538) );
  OR2X1_RVT U6535 ( .A1(n6540), .A2(n12394), .Y(n6537) );
  OR2X1_RVT U6536 ( .A1(n6542), .A2(n12385), .Y(n6531) );
  AND4X1_RVT U6537 ( .A1(n6543), .A2(n6544), .A3(n6545), .A4(n6546), .Y(n6542)
         );
  OR2X1_RVT U6538 ( .A1(n6547), .A2(n6548), .Y(n6546) );
  OR2X1_RVT U6539 ( .A1(n12402), .A2(n12397), .Y(n6548) );
  AND2X1_RVT U6540 ( .A1(n6549), .A2(n6550), .Y(n6545) );
  OR2X1_RVT U6541 ( .A1(n12802), .A2(n6551), .Y(n6544) );
  OR2X1_RVT U6542 ( .A1(n6552), .A2(n6553), .Y(n6543) );
  AND2X1_RVT U6543 ( .A1(n6554), .A2(n6555), .Y(n6552) );
  OR2X1_RVT U6544 ( .A1(n12402), .A2(n6556), .Y(n6555) );
  OR2X1_RVT U6545 ( .A1(n6489), .A2(n6557), .Y(n6530) );
  OR2X1_RVT U6546 ( .A1(n6556), .A2(n6558), .Y(n6529) );
  OR2X1_RVT U6547 ( .A1(n6559), .A2(n6560), .Y(n6527) );
  OR2X1_RVT U6548 ( .A1(n6561), .A2(n6554), .Y(n6526) );
  OR2X1_RVT U6549 ( .A1(n6562), .A2(n6563), .Y(n6525) );
  AND4X1_RVT U6550 ( .A1(n6564), .A2(n6565), .A3(n6566), .A4(n6567), .Y(n6466)
         );
  AND2X1_RVT U6551 ( .A1(n6568), .A2(n6569), .Y(n6567) );
  OR2X1_RVT U6552 ( .A1(n6553), .A2(n6570), .Y(n6569) );
  AND2X1_RVT U6553 ( .A1(n6571), .A2(n6572), .Y(n6568) );
  OR2X1_RVT U6554 ( .A1(n6573), .A2(n6496), .Y(n6572) );
  OR2X1_RVT U6555 ( .A1(n6497), .A2(n6574), .Y(n6571) );
  OR2X1_RVT U6556 ( .A1(n174), .A2(n6575), .Y(n6566) );
  OR2X1_RVT U6557 ( .A1(n6576), .A2(n12392), .Y(n6565) );
  OR2X1_RVT U6558 ( .A1(n12395), .A2(n6578), .Y(n6564) );
  AND4X1_RVT U6559 ( .A1(n6580), .A2(n6581), .A3(n6582), .A4(n6583), .Y(n6579)
         );
  AND4X1_RVT U6560 ( .A1(n6584), .A2(n6475), .A3(n6585), .A4(n6586), .Y(n6583)
         );
  AND4X1_RVT U6561 ( .A1(n6587), .A2(n6588), .A3(n6589), .A4(n6590), .Y(n6586)
         );
  OR2X1_RVT U6562 ( .A1(n6496), .A2(n6591), .Y(n6590) );
  OR2X1_RVT U6563 ( .A1(n6592), .A2(n12407), .Y(n6591) );
  OR2X1_RVT U6564 ( .A1(n6497), .A2(n6593), .Y(n6589) );
  OR2X1_RVT U6565 ( .A1(n174), .A2(n12391), .Y(n6593) );
  OR2X1_RVT U6566 ( .A1(n6594), .A2(n6540), .Y(n6588) );
  AND2X1_RVT U6567 ( .A1(n6551), .A2(n6595), .Y(n6594) );
  OR2X1_RVT U6568 ( .A1(n6596), .A2(n6597), .Y(n6587) );
  AND2X1_RVT U6569 ( .A1(n6598), .A2(n6599), .Y(n6596) );
  AND2X1_RVT U6570 ( .A1(n6600), .A2(n6601), .Y(n6585) );
  OR2X1_RVT U6571 ( .A1(n6547), .A2(n6602), .Y(n6601) );
  OR2X1_RVT U6572 ( .A1(n6603), .A2(n12800), .Y(n6602) );
  OR2X1_RVT U6573 ( .A1(n6604), .A2(n6605), .Y(n6600) );
  OR2X1_RVT U6574 ( .A1(n6606), .A2(n12396), .Y(n6605) );
  OR2X1_RVT U6575 ( .A1(n6482), .A2(n6607), .Y(n6475) );
  AND4X1_RVT U6576 ( .A1(n6608), .A2(n6609), .A3(n6610), .A4(n6611), .Y(n6582)
         );
  AND4X1_RVT U6577 ( .A1(n6612), .A2(n6613), .A3(n6614), .A4(n6615), .Y(n6611)
         );
  OR2X1_RVT U6578 ( .A1(n6616), .A2(n12410), .Y(n6615) );
  AND2X1_RVT U6579 ( .A1(n6618), .A2(n6619), .Y(n6616) );
  OR2X1_RVT U6580 ( .A1(n12379), .A2(n6497), .Y(n6619) );
  OR2X1_RVT U6581 ( .A1(n6620), .A2(n6499), .Y(n6614) );
  AND2X1_RVT U6582 ( .A1(n6621), .A2(n6622), .Y(n6620) );
  OR2X1_RVT U6583 ( .A1(n6623), .A2(n12799), .Y(n6613) );
  AND2X1_RVT U6584 ( .A1(n6624), .A2(n6625), .Y(n6623) );
  OR2X1_RVT U6585 ( .A1(n6626), .A2(n6575), .Y(n6625) );
  AND2X1_RVT U6586 ( .A1(n12410), .A2(n12394), .Y(n6626) );
  OR2X1_RVT U6587 ( .A1(n6627), .A2(n12380), .Y(n6612) );
  AND2X1_RVT U6588 ( .A1(n6629), .A2(n6630), .Y(n6627) );
  OR2X1_RVT U6589 ( .A1(n6631), .A2(n12386), .Y(n6610) );
  AND2X1_RVT U6590 ( .A1(n6632), .A2(n6633), .Y(n6631) );
  OR2X1_RVT U6591 ( .A1(n12394), .A2(n6634), .Y(n6633) );
  AND2X1_RVT U6592 ( .A1(n6635), .A2(n6636), .Y(n6632) );
  OR2X1_RVT U6593 ( .A1(n6637), .A2(n6638), .Y(n6635) );
  OR2X1_RVT U6594 ( .A1(n6482), .A2(n6553), .Y(n6638) );
  OR2X1_RVT U6595 ( .A1(n6639), .A2(n12796), .Y(n6609) );
  AND2X1_RVT U6596 ( .A1(n6640), .A2(n6641), .Y(n6639) );
  OR2X1_RVT U6597 ( .A1(n6642), .A2(n6643), .Y(n6608) );
  AND2X1_RVT U6598 ( .A1(n6644), .A2(n6645), .Y(n6642) );
  AND2X1_RVT U6599 ( .A1(n6646), .A2(n6647), .Y(n6644) );
  OR2X1_RVT U6600 ( .A1(n176), .A2(n6575), .Y(n6647) );
  OR2X1_RVT U6601 ( .A1(n12404), .A2(n6540), .Y(n6646) );
  AND4X1_RVT U6602 ( .A1(n6648), .A2(n6649), .A3(n6650), .A4(n6651), .Y(n6581)
         );
  AND4X1_RVT U6603 ( .A1(n6652), .A2(n6653), .A3(n6654), .A4(n6655), .Y(n6651)
         );
  OR2X1_RVT U6604 ( .A1(n6575), .A2(n6574), .Y(n6655) );
  OR2X1_RVT U6605 ( .A1(n6506), .A2(n6656), .Y(n6654) );
  OR2X1_RVT U6606 ( .A1(n6539), .A2(n6657), .Y(n6653) );
  OR2X1_RVT U6607 ( .A1(n6482), .A2(n6658), .Y(n6652) );
  AND2X1_RVT U6608 ( .A1(n6659), .A2(n6660), .Y(n6650) );
  OR2X1_RVT U6609 ( .A1(n12405), .A2(n6661), .Y(n6660) );
  OR2X1_RVT U6610 ( .A1(n12384), .A2(n6558), .Y(n6659) );
  OR2X1_RVT U6611 ( .A1(n6662), .A2(n6517), .Y(n6649) );
  AND4X1_RVT U6612 ( .A1(n6663), .A2(n6664), .A3(n6665), .A4(n6666), .Y(n6662)
         );
  OR2X1_RVT U6613 ( .A1(n6667), .A2(n6482), .Y(n6665) );
  OR2X1_RVT U6614 ( .A1(n12788), .A2(n6668), .Y(n6664) );
  OR2X1_RVT U6615 ( .A1(n6669), .A2(n12796), .Y(n6663) );
  AND2X1_RVT U6616 ( .A1(n6560), .A2(n6670), .Y(n6669) );
  OR2X1_RVT U6617 ( .A1(n6562), .A2(n6671), .Y(n6648) );
  AND4X1_RVT U6618 ( .A1(n6672), .A2(n6673), .A3(n6674), .A4(n6675), .Y(n6580)
         );
  AND4X1_RVT U6619 ( .A1(n6676), .A2(n6677), .A3(n6678), .A4(n6679), .Y(n6675)
         );
  OR2X1_RVT U6620 ( .A1(n12792), .A2(n6680), .Y(n6679) );
  OR2X1_RVT U6621 ( .A1(n12793), .A2(n6681), .Y(n6678) );
  OR2X1_RVT U6622 ( .A1(n12790), .A2(n6682), .Y(n6677) );
  OR2X1_RVT U6623 ( .A1(n12378), .A2(n6683), .Y(n6676) );
  OR2X1_RVT U6624 ( .A1(n6684), .A2(n12385), .Y(n6673) );
  AND4X1_RVT U6625 ( .A1(n6686), .A2(n6687), .A3(n6688), .A4(n6689), .Y(n6685)
         );
  AND4X1_RVT U6626 ( .A1(n6690), .A2(n6691), .A3(n6692), .A4(n6693), .Y(n6689)
         );
  AND4X1_RVT U6627 ( .A1(n6694), .A2(n6471), .A3(n6641), .A4(n6695), .Y(n6693)
         );
  OR2X1_RVT U6628 ( .A1(n6696), .A2(n12787), .Y(n6471) );
  AND2X1_RVT U6629 ( .A1(n6697), .A2(n6698), .Y(n6696) );
  OR2X1_RVT U6630 ( .A1(n6515), .A2(n6699), .Y(n6698) );
  OR2X1_RVT U6631 ( .A1(n6700), .A2(n6597), .Y(n6697) );
  OR2X1_RVT U6632 ( .A1(n6701), .A2(n6556), .Y(n6694) );
  AND2X1_RVT U6633 ( .A1(n6702), .A2(n6703), .Y(n6701) );
  OR2X1_RVT U6634 ( .A1(n12792), .A2(n6540), .Y(n6703) );
  OR2X1_RVT U6635 ( .A1(n6704), .A2(n6499), .Y(n6692) );
  AND2X1_RVT U6636 ( .A1(n6705), .A2(n6706), .Y(n6704) );
  OR2X1_RVT U6637 ( .A1(n6707), .A2(n12798), .Y(n6706) );
  AND2X1_RVT U6638 ( .A1(n6547), .A2(n6708), .Y(n6707) );
  OR2X1_RVT U6639 ( .A1(n6709), .A2(n12405), .Y(n6691) );
  AND2X1_RVT U6640 ( .A1(n6710), .A2(n6711), .Y(n6709) );
  OR2X1_RVT U6641 ( .A1(n6540), .A2(n6506), .Y(n6711) );
  OR2X1_RVT U6642 ( .A1(n6712), .A2(n12388), .Y(n6690) );
  AND2X1_RVT U6643 ( .A1(n6624), .A2(n6713), .Y(n6712) );
  OR2X1_RVT U6644 ( .A1(n6553), .A2(n6714), .Y(n6624) );
  AND4X1_RVT U6645 ( .A1(n6715), .A2(n6716), .A3(n6717), .A4(n6718), .Y(n6688)
         );
  OR2X1_RVT U6646 ( .A1(n6719), .A2(n12395), .Y(n6718) );
  AND2X1_RVT U6647 ( .A1(n6720), .A2(n6721), .Y(n6719) );
  OR2X1_RVT U6648 ( .A1(n6597), .A2(n6497), .Y(n6721) );
  AND2X1_RVT U6649 ( .A1(n6722), .A2(n6723), .Y(n6720) );
  OR2X1_RVT U6650 ( .A1(n6637), .A2(n6699), .Y(n6722) );
  AND2X1_RVT U6651 ( .A1(n6724), .A2(n6725), .Y(n6717) );
  OR2X1_RVT U6652 ( .A1(n6726), .A2(n6628), .Y(n6725) );
  AND2X1_RVT U6653 ( .A1(n6727), .A2(n6536), .Y(n6726) );
  OR2X1_RVT U6654 ( .A1(n6482), .A2(n6597), .Y(n6536) );
  OR2X1_RVT U6655 ( .A1(n6728), .A2(n176), .Y(n6724) );
  AND2X1_RVT U6656 ( .A1(n6729), .A2(n6730), .Y(n6728) );
  OR2X1_RVT U6657 ( .A1(n6731), .A2(n12397), .Y(n6730) );
  AND2X1_RVT U6658 ( .A1(n6732), .A2(n6733), .Y(n6731) );
  OR2X1_RVT U6659 ( .A1(n12392), .A2(n6547), .Y(n6733) );
  OR2X1_RVT U6660 ( .A1(n12802), .A2(n12394), .Y(n6732) );
  AND2X1_RVT U6661 ( .A1(n6598), .A2(n6708), .Y(n6729) );
  OR2X1_RVT U6662 ( .A1(n6628), .A2(n6734), .Y(n6598) );
  OR2X1_RVT U6663 ( .A1(n12797), .A2(n12793), .Y(n6734) );
  OR2X1_RVT U6664 ( .A1(n6735), .A2(n6617), .Y(n6716) );
  AND4X1_RVT U6665 ( .A1(n6576), .A2(n6736), .A3(n6737), .A4(n6738), .Y(n6735)
         );
  OR2X1_RVT U6666 ( .A1(n12396), .A2(n6597), .Y(n6738) );
  AND2X1_RVT U6667 ( .A1(n6739), .A2(n6740), .Y(n6737) );
  OR2X1_RVT U6668 ( .A1(n12802), .A2(n12405), .Y(n6736) );
  AND2X1_RVT U6669 ( .A1(n6741), .A2(n6742), .Y(n6576) );
  OR2X1_RVT U6670 ( .A1(n6743), .A2(n174), .Y(n6742) );
  OR2X1_RVT U6671 ( .A1(n6540), .A2(n12787), .Y(n6741) );
  AND2X1_RVT U6672 ( .A1(n6744), .A2(n6745), .Y(n6715) );
  OR2X1_RVT U6673 ( .A1(n6746), .A2(n12789), .Y(n6745) );
  AND2X1_RVT U6674 ( .A1(n6747), .A2(n6748), .Y(n6746) );
  OR2X1_RVT U6675 ( .A1(n6749), .A2(n12399), .Y(n6748) );
  AND2X1_RVT U6676 ( .A1(n6750), .A2(n6751), .Y(n6749) );
  AND2X1_RVT U6677 ( .A1(n6752), .A2(n6753), .Y(n6747) );
  OR2X1_RVT U6678 ( .A1(n6754), .A2(n12408), .Y(n6744) );
  AND4X1_RVT U6679 ( .A1(n6755), .A2(n6756), .A3(n6757), .A4(n6758), .Y(n6754)
         );
  OR2X1_RVT U6680 ( .A1(n12801), .A2(n6759), .Y(n6757) );
  OR2X1_RVT U6681 ( .A1(n174), .A2(n6554), .Y(n6756) );
  OR2X1_RVT U6682 ( .A1(n6643), .A2(n6597), .Y(n6755) );
  AND4X1_RVT U6683 ( .A1(n6760), .A2(n6761), .A3(n6762), .A4(n6763), .Y(n6687)
         );
  AND2X1_RVT U6684 ( .A1(n6764), .A2(n6607), .Y(n6763) );
  OR2X1_RVT U6685 ( .A1(n12383), .A2(n6573), .Y(n6607) );
  AND2X1_RVT U6686 ( .A1(n6765), .A2(n6766), .Y(n6764) );
  OR2X1_RVT U6687 ( .A1(n6767), .A2(n6522), .Y(n6766) );
  OR2X1_RVT U6688 ( .A1(n6574), .A2(n6634), .Y(n6765) );
  OR2X1_RVT U6689 ( .A1(n174), .A2(n6768), .Y(n6762) );
  OR2X1_RVT U6690 ( .A1(n12800), .A2(n6769), .Y(n6761) );
  OR2X1_RVT U6691 ( .A1(n6643), .A2(n6770), .Y(n6760) );
  AND4X1_RVT U6692 ( .A1(n6771), .A2(n6772), .A3(n6773), .A4(n6774), .Y(n6686)
         );
  AND2X1_RVT U6693 ( .A1(n6775), .A2(n6776), .Y(n6774) );
  OR2X1_RVT U6694 ( .A1(n12378), .A2(n6777), .Y(n6776) );
  AND2X1_RVT U6695 ( .A1(n6778), .A2(n6779), .Y(n6775) );
  OR2X1_RVT U6696 ( .A1(n6539), .A2(n6549), .Y(n6779) );
  OR2X1_RVT U6697 ( .A1(n12399), .A2(n6599), .Y(n6549) );
  OR2X1_RVT U6698 ( .A1(n12385), .A2(n6780), .Y(n6778) );
  OR2X1_RVT U6699 ( .A1(n6520), .A2(n6513), .Y(n6773) );
  OR2X1_RVT U6700 ( .A1(n6606), .A2(n6781), .Y(n6513) );
  OR2X1_RVT U6701 ( .A1(n12796), .A2(n6782), .Y(n6772) );
  OR2X1_RVT U6702 ( .A1(n12397), .A2(n6640), .Y(n6771) );
  OR2X1_RVT U6703 ( .A1(n12787), .A2(n6702), .Y(n6640) );
  AND4X1_RVT U6704 ( .A1(n6784), .A2(n6785), .A3(n6786), .A4(n6787), .Y(n6783)
         );
  AND4X1_RVT U6705 ( .A1(n6788), .A2(n6789), .A3(n6790), .A4(n6791), .Y(n6787)
         );
  OR2X1_RVT U6706 ( .A1(n184), .A2(n6792), .Y(n6791) );
  OR2X1_RVT U6707 ( .A1(n6793), .A2(n12410), .Y(n6792) );
  AND2X1_RVT U6708 ( .A1(n12399), .A2(n6559), .Y(n6793) );
  AND2X1_RVT U6709 ( .A1(n6474), .A2(n6794), .Y(n6790) );
  OR2X1_RVT U6710 ( .A1(n12388), .A2(n6795), .Y(n6474) );
  OR2X1_RVT U6711 ( .A1(n184), .A2(n6553), .Y(n6795) );
  OR2X1_RVT U6712 ( .A1(n6796), .A2(n6482), .Y(n6789) );
  AND2X1_RVT U6713 ( .A1(n6797), .A2(n6798), .Y(n6796) );
  AND2X1_RVT U6714 ( .A1(n6799), .A2(n6800), .Y(n6788) );
  OR2X1_RVT U6715 ( .A1(n6801), .A2(n6802), .Y(n6800) );
  AND2X1_RVT U6716 ( .A1(n6803), .A2(n6563), .Y(n6801) );
  OR2X1_RVT U6717 ( .A1(n6804), .A2(n6554), .Y(n6799) );
  AND2X1_RVT U6718 ( .A1(n6739), .A2(n6573), .Y(n6804) );
  OR2X1_RVT U6719 ( .A1(n12386), .A2(n6805), .Y(n6739) );
  OR2X1_RVT U6720 ( .A1(n12802), .A2(n12396), .Y(n6805) );
  AND4X1_RVT U6721 ( .A1(n6806), .A2(n6807), .A3(n6808), .A4(n6809), .Y(n6786)
         );
  OR2X1_RVT U6722 ( .A1(n6810), .A2(n12792), .Y(n6809) );
  AND2X1_RVT U6723 ( .A1(n6622), .A2(n6811), .Y(n6810) );
  OR2X1_RVT U6724 ( .A1(n12800), .A2(n6667), .Y(n6622) );
  AND2X1_RVT U6725 ( .A1(n6812), .A2(n6813), .Y(n6808) );
  OR2X1_RVT U6726 ( .A1(n6814), .A2(n12790), .Y(n6813) );
  AND2X1_RVT U6727 ( .A1(n6815), .A2(n6816), .Y(n6814) );
  OR2X1_RVT U6728 ( .A1(n6517), .A2(n6759), .Y(n6816) );
  OR2X1_RVT U6729 ( .A1(n6817), .A2(n12788), .Y(n6812) );
  AND2X1_RVT U6730 ( .A1(n6818), .A2(n6819), .Y(n6817) );
  OR2X1_RVT U6731 ( .A1(n6820), .A2(n12399), .Y(n6807) );
  AND2X1_RVT U6732 ( .A1(n6821), .A2(n6822), .Y(n6820) );
  AND2X1_RVT U6733 ( .A1(n6823), .A2(n6824), .Y(n6821) );
  AND2X1_RVT U6734 ( .A1(n6825), .A2(n6826), .Y(n6806) );
  OR2X1_RVT U6735 ( .A1(n6827), .A2(n6743), .Y(n6826) );
  AND2X1_RVT U6736 ( .A1(n6828), .A2(n6574), .Y(n6827) );
  AND2X1_RVT U6737 ( .A1(n6829), .A2(n6830), .Y(n6828) );
  OR2X1_RVT U6738 ( .A1(n6831), .A2(n12402), .Y(n6825) );
  AND2X1_RVT U6739 ( .A1(n6832), .A2(n6833), .Y(n6831) );
  OR2X1_RVT U6740 ( .A1(n12799), .A2(n12404), .Y(n6833) );
  AND2X1_RVT U6741 ( .A1(n6563), .A2(n6834), .Y(n6832) );
  AND4X1_RVT U6742 ( .A1(n6835), .A2(n6836), .A3(n6837), .A4(n6838), .Y(n6785)
         );
  AND2X1_RVT U6743 ( .A1(n6839), .A2(n6840), .Y(n6838) );
  OR2X1_RVT U6744 ( .A1(n6556), .A2(n6630), .Y(n6840) );
  OR2X1_RVT U6745 ( .A1(n12794), .A2(n6563), .Y(n6630) );
  AND2X1_RVT U6746 ( .A1(n6841), .A2(n6842), .Y(n6839) );
  OR2X1_RVT U6747 ( .A1(n6708), .A2(n6522), .Y(n6842) );
  OR2X1_RVT U6748 ( .A1(n12801), .A2(n12395), .Y(n6522) );
  OR2X1_RVT U6749 ( .A1(n6606), .A2(n6656), .Y(n6841) );
  OR2X1_RVT U6750 ( .A1(n12789), .A2(n6843), .Y(n6656) );
  OR2X1_RVT U6751 ( .A1(n6844), .A2(n12378), .Y(n6837) );
  AND4X1_RVT U6752 ( .A1(n6845), .A2(n6846), .A3(n6847), .A4(n6848), .Y(n6844)
         );
  OR2X1_RVT U6753 ( .A1(n6781), .A2(n6554), .Y(n6847) );
  OR2X1_RVT U6754 ( .A1(n6849), .A2(n6551), .Y(n6846) );
  OR2X1_RVT U6755 ( .A1(n12798), .A2(n6506), .Y(n6845) );
  OR2X1_RVT U6756 ( .A1(n6850), .A2(n12379), .Y(n6836) );
  AND2X1_RVT U6757 ( .A1(n6851), .A2(n6852), .Y(n6850) );
  OR2X1_RVT U6758 ( .A1(n6781), .A2(n6506), .Y(n6852) );
  AND2X1_RVT U6759 ( .A1(n6853), .A2(n6782), .Y(n6851) );
  OR2X1_RVT U6760 ( .A1(n6554), .A2(n6854), .Y(n6782) );
  OR2X1_RVT U6761 ( .A1(n12789), .A2(n12801), .Y(n6854) );
  OR2X1_RVT U6762 ( .A1(n6855), .A2(n12386), .Y(n6835) );
  AND4X1_RVT U6763 ( .A1(n6856), .A2(n6769), .A3(n6578), .A4(n6550), .Y(n6855)
         );
  OR2X1_RVT U6764 ( .A1(n6575), .A2(n6857), .Y(n6550) );
  OR2X1_RVT U6765 ( .A1(n12791), .A2(n6512), .Y(n6857) );
  OR2X1_RVT U6766 ( .A1(n6637), .A2(n6671), .Y(n6578) );
  OR2X1_RVT U6767 ( .A1(n6556), .A2(n6858), .Y(n6769) );
  OR2X1_RVT U6768 ( .A1(n12410), .A2(n12379), .Y(n6858) );
  OR2X1_RVT U6769 ( .A1(n6515), .A2(n6859), .Y(n6856) );
  OR2X1_RVT U6770 ( .A1(n6860), .A2(n12384), .Y(n6859) );
  AND4X1_RVT U6771 ( .A1(n6861), .A2(n6862), .A3(n6863), .A4(n6864), .Y(n6784)
         );
  AND2X1_RVT U6772 ( .A1(n6865), .A2(n6866), .Y(n6864) );
  AND2X1_RVT U6773 ( .A1(n6867), .A2(n6868), .Y(n6865) );
  OR2X1_RVT U6774 ( .A1(n6547), .A2(n6822), .Y(n6868) );
  OR2X1_RVT U6775 ( .A1(n6559), .A2(n6869), .Y(n6822) );
  OR2X1_RVT U6776 ( .A1(n12790), .A2(n12792), .Y(n6869) );
  OR2X1_RVT U6777 ( .A1(n12797), .A2(n6870), .Y(n6867) );
  OR2X1_RVT U6778 ( .A1(n12395), .A2(n6871), .Y(n6863) );
  OR2X1_RVT U6779 ( .A1(n12800), .A2(n6872), .Y(n6862) );
  OR2X1_RVT U6780 ( .A1(n6559), .A2(n6873), .Y(n6861) );
  AND4X1_RVT U6781 ( .A1(n6875), .A2(n6876), .A3(n6877), .A4(n6878), .Y(n6874)
         );
  AND4X1_RVT U6782 ( .A1(n6879), .A2(n6880), .A3(n6881), .A4(n6882), .Y(n6878)
         );
  AND4X1_RVT U6783 ( .A1(n6883), .A2(n6884), .A3(n6476), .A4(n6885), .Y(n6882)
         );
  OR2X1_RVT U6784 ( .A1(n6617), .A2(n6886), .Y(n6476) );
  OR2X1_RVT U6785 ( .A1(n6708), .A2(n176), .Y(n6886) );
  OR2X1_RVT U6786 ( .A1(n6480), .A2(n6887), .Y(n6884) );
  OR2X1_RVT U6787 ( .A1(n12795), .A2(n12798), .Y(n6887) );
  OR2X1_RVT U6788 ( .A1(n6743), .A2(n6888), .Y(n6883) );
  OR2X1_RVT U6789 ( .A1(n6889), .A2(n6517), .Y(n6888) );
  AND2X1_RVT U6790 ( .A1(n12399), .A2(n6617), .Y(n6889) );
  OR2X1_RVT U6791 ( .A1(n6890), .A2(n12405), .Y(n6881) );
  AND2X1_RVT U6792 ( .A1(n6758), .A2(n6830), .Y(n6890) );
  OR2X1_RVT U6793 ( .A1(n176), .A2(n6891), .Y(n6830) );
  OR2X1_RVT U6794 ( .A1(n12378), .A2(n12794), .Y(n6891) );
  OR2X1_RVT U6795 ( .A1(n6547), .A2(n6892), .Y(n6758) );
  OR2X1_RVT U6796 ( .A1(n12792), .A2(n6539), .Y(n6892) );
  OR2X1_RVT U6797 ( .A1(n6893), .A2(n6497), .Y(n6880) );
  AND2X1_RVT U6798 ( .A1(n6894), .A2(n6702), .Y(n6893) );
  OR2X1_RVT U6799 ( .A1(n6603), .A2(n6597), .Y(n6879) );
  AND4X1_RVT U6800 ( .A1(n6895), .A2(n6896), .A3(n6897), .A4(n6898), .Y(n6877)
         );
  AND2X1_RVT U6801 ( .A1(n6899), .A2(n6900), .Y(n6898) );
  OR2X1_RVT U6802 ( .A1(n6901), .A2(n12399), .Y(n6900) );
  AND2X1_RVT U6803 ( .A1(n6902), .A2(n6570), .Y(n6901) );
  AND2X1_RVT U6804 ( .A1(n6903), .A2(n6904), .Y(n6899) );
  OR2X1_RVT U6805 ( .A1(n6905), .A2(n6553), .Y(n6904) );
  AND2X1_RVT U6806 ( .A1(n6524), .A2(n6496), .Y(n6905) );
  OR2X1_RVT U6807 ( .A1(n12800), .A2(n6595), .Y(n6524) );
  OR2X1_RVT U6808 ( .A1(n6906), .A2(n6606), .Y(n6903) );
  AND2X1_RVT U6809 ( .A1(n6798), .A2(n6907), .Y(n6906) );
  OR2X1_RVT U6810 ( .A1(n12801), .A2(n6634), .Y(n6798) );
  OR2X1_RVT U6811 ( .A1(n6908), .A2(n12792), .Y(n6897) );
  AND2X1_RVT U6812 ( .A1(n6501), .A2(n6909), .Y(n6908) );
  OR2X1_RVT U6813 ( .A1(n6637), .A2(n6561), .Y(n6909) );
  OR2X1_RVT U6814 ( .A1(n6540), .A2(n6743), .Y(n6501) );
  OR2X1_RVT U6815 ( .A1(n6910), .A2(n174), .Y(n6896) );
  AND2X1_RVT U6816 ( .A1(n6551), .A2(n6911), .Y(n6910) );
  OR2X1_RVT U6817 ( .A1(n6912), .A2(n12383), .Y(n6911) );
  AND2X1_RVT U6818 ( .A1(n6913), .A2(n6914), .Y(n6912) );
  OR2X1_RVT U6819 ( .A1(n12793), .A2(n6534), .Y(n6914) );
  OR2X1_RVT U6820 ( .A1(n12410), .A2(n6637), .Y(n6551) );
  OR2X1_RVT U6821 ( .A1(n6915), .A2(n6621), .Y(n6895) );
  AND2X1_RVT U6822 ( .A1(n6554), .A2(n6599), .Y(n6915) );
  OR2X1_RVT U6823 ( .A1(n12789), .A2(n6482), .Y(n6599) );
  AND4X1_RVT U6824 ( .A1(n6916), .A2(n6917), .A3(n6918), .A4(n6919), .Y(n6876)
         );
  AND4X1_RVT U6825 ( .A1(n6920), .A2(n6921), .A3(n6922), .A4(n6923), .Y(n6919)
         );
  OR2X1_RVT U6826 ( .A1(n6924), .A2(n12800), .Y(n6923) );
  AND2X1_RVT U6827 ( .A1(n6657), .A2(n6925), .Y(n6924) );
  OR2X1_RVT U6828 ( .A1(n12407), .A2(n6506), .Y(n6925) );
  OR2X1_RVT U6829 ( .A1(n6926), .A2(n6499), .Y(n6922) );
  AND2X1_RVT U6830 ( .A1(n6927), .A2(n6928), .Y(n6926) );
  OR2X1_RVT U6831 ( .A1(n6929), .A2(n6534), .Y(n6928) );
  AND2X1_RVT U6832 ( .A1(n6559), .A2(n6547), .Y(n6929) );
  AND2X1_RVT U6833 ( .A1(n6561), .A2(n6803), .Y(n6927) );
  OR2X1_RVT U6834 ( .A1(n12408), .A2(n6699), .Y(n6803) );
  OR2X1_RVT U6835 ( .A1(n6930), .A2(n12397), .Y(n6921) );
  AND2X1_RVT U6836 ( .A1(n6931), .A2(n6932), .Y(n6930) );
  OR2X1_RVT U6837 ( .A1(n6547), .A2(n6933), .Y(n6932) );
  AND2X1_RVT U6838 ( .A1(n6629), .A2(n6823), .Y(n6931) );
  OR2X1_RVT U6839 ( .A1(n6539), .A2(n6714), .Y(n6823) );
  OR2X1_RVT U6840 ( .A1(n6512), .A2(n6934), .Y(n6629) );
  OR2X1_RVT U6841 ( .A1(n6935), .A2(n6482), .Y(n6920) );
  AND4X1_RVT U6842 ( .A1(n6936), .A2(n6937), .A3(n6938), .A4(n6871), .Y(n6935)
         );
  OR2X1_RVT U6843 ( .A1(n6575), .A2(n6939), .Y(n6871) );
  OR2X1_RVT U6844 ( .A1(n12378), .A2(n6539), .Y(n6939) );
  OR2X1_RVT U6845 ( .A1(n12797), .A2(n6781), .Y(n6937) );
  OR2X1_RVT U6846 ( .A1(n6540), .A2(n6637), .Y(n6936) );
  OR2X1_RVT U6847 ( .A1(n6708), .A2(n6750), .Y(n6918) );
  OR2X1_RVT U6848 ( .A1(n6940), .A2(n12381), .Y(n6917) );
  AND4X1_RVT U6849 ( .A1(n6941), .A2(n6942), .A3(n6584), .A4(n6682), .Y(n6940)
         );
  OR2X1_RVT U6850 ( .A1(n6506), .A2(n6671), .Y(n6682) );
  OR2X1_RVT U6851 ( .A1(n12797), .A2(n174), .Y(n6671) );
  OR2X1_RVT U6852 ( .A1(n6499), .A2(n6563), .Y(n6584) );
  OR2X1_RVT U6853 ( .A1(n12789), .A2(n6934), .Y(n6916) );
  AND4X1_RVT U6854 ( .A1(n6943), .A2(n6944), .A3(n6945), .A4(n6946), .Y(n6875)
         );
  OR2X1_RVT U6855 ( .A1(n12386), .A2(n6947), .Y(n6946) );
  AND2X1_RVT U6856 ( .A1(n6948), .A2(n6949), .Y(n6945) );
  OR2X1_RVT U6857 ( .A1(n12407), .A2(n6702), .Y(n6949) );
  OR2X1_RVT U6858 ( .A1(n6489), .A2(n6563), .Y(n6948) );
  OR2X1_RVT U6859 ( .A1(n176), .A2(n6520), .Y(n6563) );
  OR2X1_RVT U6860 ( .A1(n12410), .A2(n6681), .Y(n6944) );
  OR2X1_RVT U6861 ( .A1(n6556), .A2(n6950), .Y(n6681) );
  AND2X1_RVT U6862 ( .A1(n6951), .A2(n6952), .Y(n6943) );
  OR2X1_RVT U6863 ( .A1(n12379), .A2(n6953), .Y(n6952) );
  OR2X1_RVT U6864 ( .A1(n6559), .A2(n6508), .Y(n6951) );
  OR2X1_RVT U6865 ( .A1(n6482), .A2(n6767), .Y(n6508) );
  AND4X1_RVT U6866 ( .A1(n6955), .A2(n6956), .A3(n6957), .A4(n6958), .Y(n6954)
         );
  AND4X1_RVT U6867 ( .A1(n6959), .A2(n6960), .A3(n6961), .A4(n6962), .Y(n6958)
         );
  AND4X1_RVT U6868 ( .A1(n6963), .A2(n6964), .A3(n6123), .A4(n6965), .Y(n6962)
         );
  OR2X1_RVT U6869 ( .A1(n1332), .A2(n6191), .Y(n6123) );
  AND2X1_RVT U6870 ( .A1(n6966), .A2(n6967), .Y(n6961) );
  OR2X1_RVT U6871 ( .A1(n1323), .A2(n6968), .Y(n6966) );
  OR2X1_RVT U6872 ( .A1(n12872), .A2(n12190), .Y(n6968) );
  OR2X1_RVT U6873 ( .A1(n6969), .A2(n12206), .Y(n6960) );
  AND2X1_RVT U6874 ( .A1(n1313), .A2(n6970), .Y(n6969) );
  OR2X1_RVT U6875 ( .A1(n6971), .A2(n12209), .Y(n6970) );
  AND2X1_RVT U6876 ( .A1(n6972), .A2(n6973), .Y(n6971) );
  OR2X1_RVT U6877 ( .A1(n6974), .A2(n12212), .Y(n6959) );
  AND2X1_RVT U6878 ( .A1(n6975), .A2(n6976), .Y(n6974) );
  AND4X1_RVT U6879 ( .A1(n6977), .A2(n6978), .A3(n6979), .A4(n6980), .Y(n6957)
         );
  AND4X1_RVT U6880 ( .A1(n6981), .A2(n6982), .A3(n6983), .A4(n6984), .Y(n6980)
         );
  OR2X1_RVT U6881 ( .A1(n6985), .A2(n85), .Y(n6984) );
  AND2X1_RVT U6882 ( .A1(n6986), .A2(n6987), .Y(n6985) );
  OR2X1_RVT U6883 ( .A1(n6988), .A2(n12149), .Y(n6987) );
  AND2X1_RVT U6884 ( .A1(n1348), .A2(n6989), .Y(n6988) );
  OR2X1_RVT U6885 ( .A1(n6990), .A2(n12195), .Y(n6983) );
  AND2X1_RVT U6886 ( .A1(n6991), .A2(n6992), .Y(n6990) );
  OR2X1_RVT U6887 ( .A1(n12876), .A2(n1359), .Y(n6992) );
  OR2X1_RVT U6888 ( .A1(n6993), .A2(n1391), .Y(n6991) );
  AND2X1_RVT U6889 ( .A1(n72), .A2(n6994), .Y(n6993) );
  OR2X1_RVT U6890 ( .A1(n12871), .A2(n12875), .Y(n6994) );
  OR2X1_RVT U6891 ( .A1(n6995), .A2(n6132), .Y(n6982) );
  AND2X1_RVT U6892 ( .A1(n6996), .A2(n6997), .Y(n6995) );
  OR2X1_RVT U6893 ( .A1(n12872), .A2(n1365), .Y(n6997) );
  AND2X1_RVT U6894 ( .A1(n6998), .A2(n6199), .Y(n6996) );
  OR2X1_RVT U6895 ( .A1(n6999), .A2(n7000), .Y(n6998) );
  OR2X1_RVT U6896 ( .A1(n7001), .A2(n12869), .Y(n6981) );
  AND2X1_RVT U6897 ( .A1(n7002), .A2(n7003), .Y(n7001) );
  OR2X1_RVT U6898 ( .A1(n76), .A2(n12206), .Y(n7003) );
  AND2X1_RVT U6899 ( .A1(n7004), .A2(n7005), .Y(n7002) );
  OR2X1_RVT U6900 ( .A1(n78), .A2(n7006), .Y(n7004) );
  OR2X1_RVT U6901 ( .A1(n7007), .A2(n7008), .Y(n6979) );
  OR2X1_RVT U6902 ( .A1(n7009), .A2(n12188), .Y(n6978) );
  AND2X1_RVT U6903 ( .A1(n7010), .A2(n7011), .Y(n7009) );
  OR2X1_RVT U6904 ( .A1(n7012), .A2(n7013), .Y(n7011) );
  AND2X1_RVT U6905 ( .A1(n7014), .A2(n7015), .Y(n7010) );
  OR2X1_RVT U6906 ( .A1(n7016), .A2(n83), .Y(n6977) );
  AND4X1_RVT U6907 ( .A1(n7017), .A2(n7018), .A3(n7019), .A4(n6196), .Y(n7016)
         );
  OR2X1_RVT U6908 ( .A1(n1314), .A2(n7000), .Y(n7018) );
  OR2X1_RVT U6909 ( .A1(n7020), .A2(n1325), .Y(n7017) );
  AND2X1_RVT U6910 ( .A1(n12195), .A2(n7021), .Y(n7020) );
  OR2X1_RVT U6911 ( .A1(n12877), .A2(n12185), .Y(n7021) );
  AND4X1_RVT U6912 ( .A1(n7022), .A2(n7023), .A3(n7024), .A4(n7025), .Y(n6956)
         );
  AND4X1_RVT U6913 ( .A1(n7026), .A2(n7027), .A3(n7028), .A4(n7029), .Y(n7025)
         );
  OR2X1_RVT U6914 ( .A1(n6197), .A2(n12926), .Y(n7029) );
  OR2X1_RVT U6915 ( .A1(n6198), .A2(n1392), .Y(n7028) );
  OR2X1_RVT U6916 ( .A1(n73), .A2(n7030), .Y(n1392) );
  OR2X1_RVT U6917 ( .A1(n1312), .A2(n7031), .Y(n7027) );
  OR2X1_RVT U6918 ( .A1(n1350), .A2(n7032), .Y(n7026) );
  OR2X1_RVT U6919 ( .A1(n12204), .A2(n7033), .Y(n7024) );
  OR2X1_RVT U6920 ( .A1(n12184), .A2(n6146), .Y(n7023) );
  OR2X1_RVT U6921 ( .A1(n12192), .A2(n1348), .Y(n6146) );
  OR2X1_RVT U6922 ( .A1(n7034), .A2(n1400), .Y(n7022) );
  AND4X1_RVT U6923 ( .A1(n7035), .A2(n7036), .A3(n1394), .A4(n7037), .Y(n6955)
         );
  AND4X1_RVT U6924 ( .A1(n7038), .A2(n7039), .A3(n7040), .A4(n7041), .Y(n7037)
         );
  OR2X1_RVT U6925 ( .A1(n12186), .A2(n7042), .Y(n7041) );
  OR2X1_RVT U6926 ( .A1(n1325), .A2(n7043), .Y(n7040) );
  OR2X1_RVT U6927 ( .A1(n12876), .A2(n7044), .Y(n7039) );
  OR2X1_RVT U6928 ( .A1(n12199), .A2(n7045), .Y(n7038) );
  AND2X1_RVT U6929 ( .A1(n7046), .A2(n7047), .Y(n1394) );
  OR2X1_RVT U6930 ( .A1(n12869), .A2(n6200), .Y(n7047) );
  OR2X1_RVT U6931 ( .A1(n7048), .A2(n83), .Y(n7046) );
  OR2X1_RVT U6932 ( .A1(n71), .A2(n7049), .Y(n7036) );
  OR2X1_RVT U6933 ( .A1(n1351), .A2(n12874), .Y(n7035) );
  AND2X1_RVT U6934 ( .A1(n7050), .A2(n7051), .Y(n1351) );
  OR2X1_RVT U6935 ( .A1(n1370), .A2(n7034), .Y(n7051) );
  OR2X1_RVT U6936 ( .A1(n7052), .A2(n12211), .Y(n7050) );
  AND4X1_RVT U6937 ( .A1(n7054), .A2(n7055), .A3(n7056), .A4(n7057), .Y(n7053)
         );
  AND4X1_RVT U6938 ( .A1(n7058), .A2(n7059), .A3(n7060), .A4(n7061), .Y(n7057)
         );
  AND4X1_RVT U6939 ( .A1(n6695), .A2(n6885), .A3(n7062), .A4(n7063), .Y(n7061)
         );
  OR2X1_RVT U6940 ( .A1(n7064), .A2(n7065), .Y(n6885) );
  OR2X1_RVT U6941 ( .A1(n6480), .A2(n6750), .Y(n6695) );
  OR2X1_RVT U6942 ( .A1(n12798), .A2(n12395), .Y(n6750) );
  AND4X1_RVT U6943 ( .A1(n6953), .A2(n6819), .A3(n6942), .A4(n6477), .Y(n7060)
         );
  OR2X1_RVT U6944 ( .A1(n7066), .A2(n6667), .Y(n6477) );
  OR2X1_RVT U6945 ( .A1(n6482), .A2(n7067), .Y(n6942) );
  OR2X1_RVT U6946 ( .A1(n6515), .A2(n174), .Y(n6819) );
  OR2X1_RVT U6947 ( .A1(n6506), .A2(n7068), .Y(n6953) );
  OR2X1_RVT U6948 ( .A1(n12385), .A2(n12405), .Y(n7068) );
  AND4X1_RVT U6949 ( .A1(n7069), .A2(n7070), .A3(n7071), .A4(n7072), .Y(n7059)
         );
  OR2X1_RVT U6950 ( .A1(n6759), .A2(n7073), .Y(n7072) );
  OR2X1_RVT U6951 ( .A1(n12405), .A2(n6539), .Y(n7073) );
  OR2X1_RVT U6952 ( .A1(n6668), .A2(n7074), .Y(n7071) );
  OR2X1_RVT U6953 ( .A1(n12799), .A2(n6556), .Y(n7074) );
  OR2X1_RVT U6954 ( .A1(n6894), .A2(n7075), .Y(n7070) );
  OR2X1_RVT U6955 ( .A1(n7076), .A2(n6553), .Y(n7075) );
  OR2X1_RVT U6956 ( .A1(n12402), .A2(n7077), .Y(n7069) );
  OR2X1_RVT U6957 ( .A1(n7078), .A2(n12385), .Y(n7077) );
  AND2X1_RVT U6958 ( .A1(n6767), .A2(n7079), .Y(n7078) );
  AND2X1_RVT U6959 ( .A1(n7080), .A2(n7081), .Y(n7058) );
  OR2X1_RVT U6960 ( .A1(n7082), .A2(n6534), .Y(n7081) );
  AND2X1_RVT U6961 ( .A1(n7083), .A2(n7084), .Y(n7082) );
  OR2X1_RVT U6962 ( .A1(n12384), .A2(n6727), .Y(n7084) );
  OR2X1_RVT U6963 ( .A1(n12388), .A2(n6802), .Y(n7083) );
  AND2X1_RVT U6964 ( .A1(n7085), .A2(n7086), .Y(n7080) );
  OR2X1_RVT U6965 ( .A1(n7087), .A2(n6573), .Y(n7086) );
  AND2X1_RVT U6966 ( .A1(n7088), .A2(n7089), .Y(n7087) );
  OR2X1_RVT U6967 ( .A1(n12391), .A2(n184), .Y(n7089) );
  NAND2X1_RVT U6968 ( .A1(n6556), .A2(n12791), .Y(n7088) );
  OR2X1_RVT U6969 ( .A1(n7090), .A2(n176), .Y(n7085) );
  AND2X1_RVT U6970 ( .A1(n6780), .A2(n6657), .Y(n7090) );
  OR2X1_RVT U6971 ( .A1(n6506), .A2(n7091), .Y(n6657) );
  OR2X1_RVT U6972 ( .A1(n12802), .A2(n12380), .Y(n7091) );
  AND4X1_RVT U6973 ( .A1(n6674), .A2(n7092), .A3(n6866), .A4(n7093), .Y(n7056)
         );
  AND4X1_RVT U6974 ( .A1(n7094), .A2(n7095), .A3(n7096), .A4(n7097), .Y(n7093)
         );
  OR2X1_RVT U6975 ( .A1(n6637), .A2(n6558), .Y(n7097) );
  OR2X1_RVT U6976 ( .A1(n6575), .A2(n6604), .Y(n7096) );
  OR2X1_RVT U6977 ( .A1(n12790), .A2(n6829), .Y(n7095) );
  OR2X1_RVT U6978 ( .A1(n6553), .A2(n6535), .Y(n6829) );
  OR2X1_RVT U6979 ( .A1(n12798), .A2(n6617), .Y(n6535) );
  OR2X1_RVT U6980 ( .A1(n12394), .A2(n6658), .Y(n7094) );
  OR2X1_RVT U6981 ( .A1(n6539), .A2(n6767), .Y(n6658) );
  OR2X1_RVT U6982 ( .A1(n12378), .A2(n6743), .Y(n6767) );
  AND2X1_RVT U6983 ( .A1(n7098), .A2(n7099), .Y(n6866) );
  OR2X1_RVT U6984 ( .A1(n7100), .A2(n6606), .Y(n7099) );
  OR2X1_RVT U6985 ( .A1(n12404), .A2(n176), .Y(n7100) );
  OR2X1_RVT U6986 ( .A1(n7101), .A2(n6489), .Y(n7098) );
  OR2X1_RVT U6987 ( .A1(n12789), .A2(n6606), .Y(n6489) );
  OR2X1_RVT U6988 ( .A1(n6503), .A2(n6553), .Y(n7101) );
  OR2X1_RVT U6989 ( .A1(n12386), .A2(n6872), .Y(n7092) );
  AND2X1_RVT U6990 ( .A1(n7102), .A2(n7103), .Y(n6674) );
  OR2X1_RVT U6991 ( .A1(n6557), .A2(n6595), .Y(n7103) );
  OR2X1_RVT U6992 ( .A1(n7104), .A2(n7105), .Y(n7102) );
  AND4X1_RVT U6993 ( .A1(n7106), .A2(n7107), .A3(n7108), .A4(n7109), .Y(n7055)
         );
  OR2X1_RVT U6994 ( .A1(n7110), .A2(n6743), .Y(n7109) );
  AND2X1_RVT U6995 ( .A1(n7111), .A2(n6752), .Y(n7110) );
  OR2X1_RVT U6996 ( .A1(n12392), .A2(n7067), .Y(n6752) );
  OR2X1_RVT U6997 ( .A1(n7112), .A2(n12795), .Y(n7108) );
  AND2X1_RVT U6998 ( .A1(n6680), .A2(n6645), .Y(n7112) );
  OR2X1_RVT U6999 ( .A1(n12789), .A2(n6621), .Y(n6645) );
  OR2X1_RVT U7000 ( .A1(n7113), .A2(n6700), .Y(n7107) );
  AND2X1_RVT U7001 ( .A1(n7114), .A2(n7115), .Y(n7113) );
  OR2X1_RVT U7002 ( .A1(n12381), .A2(n6559), .Y(n7115) );
  AND2X1_RVT U7003 ( .A1(n7116), .A2(n6597), .Y(n7114) );
  OR2X1_RVT U7004 ( .A1(n174), .A2(n6556), .Y(n7116) );
  OR2X1_RVT U7005 ( .A1(n7117), .A2(n6497), .Y(n7106) );
  AND2X1_RVT U7006 ( .A1(n7118), .A2(n7119), .Y(n7117) );
  NAND2X1_RVT U7007 ( .A1(n6482), .A2(n6860), .Y(n7119) );
  AND2X1_RVT U7008 ( .A1(n7120), .A2(n6710), .Y(n7118) );
  OR2X1_RVT U7009 ( .A1(n6643), .A2(n7067), .Y(n6710) );
  OR2X1_RVT U7010 ( .A1(n12401), .A2(n7121), .Y(n7120) );
  AND4X1_RVT U7011 ( .A1(n7122), .A2(n7123), .A3(n7124), .A4(n7125), .Y(n7054)
         );
  OR2X1_RVT U7012 ( .A1(n7126), .A2(n6520), .Y(n7125) );
  AND2X1_RVT U7013 ( .A1(n7127), .A2(n6661), .Y(n7126) );
  AND2X1_RVT U7014 ( .A1(n7128), .A2(n6683), .Y(n7127) );
  OR2X1_RVT U7015 ( .A1(n176), .A2(n7105), .Y(n6683) );
  OR2X1_RVT U7016 ( .A1(n12380), .A2(n6617), .Y(n7105) );
  OR2X1_RVT U7017 ( .A1(n7129), .A2(n12397), .Y(n7124) );
  AND2X1_RVT U7018 ( .A1(n7130), .A2(n7131), .Y(n7129) );
  OR2X1_RVT U7019 ( .A1(n7132), .A2(n12787), .Y(n7131) );
  AND2X1_RVT U7020 ( .A1(n7133), .A2(n7134), .Y(n7132) );
  OR2X1_RVT U7021 ( .A1(n12379), .A2(n6894), .Y(n7134) );
  OR2X1_RVT U7022 ( .A1(n12794), .A2(n6540), .Y(n7133) );
  AND2X1_RVT U7023 ( .A1(n7135), .A2(n7136), .Y(n7130) );
  OR2X1_RVT U7024 ( .A1(n6506), .A2(n7137), .Y(n7135) );
  OR2X1_RVT U7025 ( .A1(n7138), .A2(n6540), .Y(n7123) );
  AND4X1_RVT U7026 ( .A1(n7139), .A2(n7140), .A3(n7141), .A4(n6506), .Y(n7138)
         );
  OR2X1_RVT U7027 ( .A1(n12795), .A2(n6556), .Y(n7141) );
  OR2X1_RVT U7028 ( .A1(n12391), .A2(n6575), .Y(n7140) );
  OR2X1_RVT U7029 ( .A1(n6628), .A2(n6606), .Y(n7139) );
  OR2X1_RVT U7030 ( .A1(n7142), .A2(n6482), .Y(n7122) );
  AND4X1_RVT U7031 ( .A1(n6907), .A2(n7143), .A3(n6705), .A4(n6621), .Y(n7142)
         );
  OR2X1_RVT U7032 ( .A1(n6575), .A2(n7137), .Y(n6705) );
  OR2X1_RVT U7033 ( .A1(n6743), .A2(n6950), .Y(n7143) );
  OR2X1_RVT U7034 ( .A1(n12385), .A2(n6708), .Y(n6907) );
  AND4X1_RVT U7035 ( .A1(n7145), .A2(n7146), .A3(n7147), .A4(n7148), .Y(n7144)
         );
  AND4X1_RVT U7036 ( .A1(n6558), .A2(n6794), .A3(n7149), .A4(n7150), .Y(n7148)
         );
  AND4X1_RVT U7037 ( .A1(n6873), .A2(n6818), .A3(n7062), .A4(n7063), .Y(n7150)
         );
  OR2X1_RVT U7038 ( .A1(n7065), .A2(n6479), .Y(n7063) );
  OR2X1_RVT U7039 ( .A1(n12793), .A2(n6597), .Y(n6479) );
  OR2X1_RVT U7040 ( .A1(n6496), .A2(n7104), .Y(n7062) );
  OR2X1_RVT U7041 ( .A1(n12798), .A2(n12399), .Y(n7104) );
  OR2X1_RVT U7042 ( .A1(n12787), .A2(n6617), .Y(n6496) );
  OR2X1_RVT U7043 ( .A1(n12799), .A2(n6515), .Y(n6818) );
  OR2X1_RVT U7044 ( .A1(n12408), .A2(n12392), .Y(n6515) );
  OR2X1_RVT U7045 ( .A1(n6637), .A2(n7151), .Y(n6873) );
  OR2X1_RVT U7046 ( .A1(n12399), .A2(n6541), .Y(n7151) );
  OR2X1_RVT U7047 ( .A1(n6539), .A2(n7152), .Y(n7149) );
  OR2X1_RVT U7048 ( .A1(n6667), .A2(n12390), .Y(n7152) );
  OR2X1_RVT U7049 ( .A1(n6606), .A2(n7153), .Y(n6794) );
  OR2X1_RVT U7050 ( .A1(n6540), .A2(n12397), .Y(n7153) );
  OR2X1_RVT U7051 ( .A1(n12791), .A2(n7064), .Y(n6558) );
  OR2X1_RVT U7052 ( .A1(n12392), .A2(n6557), .Y(n7064) );
  AND4X1_RVT U7053 ( .A1(n7154), .A2(n7155), .A3(n7156), .A4(n7157), .Y(n7147)
         );
  AND4X1_RVT U7054 ( .A1(n7158), .A2(n7159), .A3(n7160), .A4(n7161), .Y(n7157)
         );
  OR2X1_RVT U7055 ( .A1(n6573), .A2(n7162), .Y(n7161) );
  OR2X1_RVT U7056 ( .A1(n12381), .A2(n6643), .Y(n7162) );
  OR2X1_RVT U7057 ( .A1(n6556), .A2(n7163), .Y(n7160) );
  OR2X1_RVT U7058 ( .A1(n7164), .A2(n6520), .Y(n7163) );
  AND2X1_RVT U7059 ( .A1(n6499), .A2(n6559), .Y(n7164) );
  OR2X1_RVT U7060 ( .A1(n7165), .A2(n7166), .Y(n7159) );
  AND2X1_RVT U7061 ( .A1(n6714), .A2(n6670), .Y(n7165) );
  OR2X1_RVT U7062 ( .A1(n12792), .A2(n184), .Y(n6670) );
  OR2X1_RVT U7063 ( .A1(n12788), .A2(n12402), .Y(n6714) );
  OR2X1_RVT U7064 ( .A1(n7167), .A2(n6554), .Y(n7158) );
  AND2X1_RVT U7065 ( .A1(n6950), .A2(n7168), .Y(n7167) );
  OR2X1_RVT U7066 ( .A1(n12790), .A2(n176), .Y(n7168) );
  OR2X1_RVT U7067 ( .A1(n7169), .A2(n12404), .Y(n7156) );
  AND2X1_RVT U7068 ( .A1(n6941), .A2(n7170), .Y(n7169) );
  OR2X1_RVT U7069 ( .A1(n6547), .A2(n6894), .Y(n7170) );
  OR2X1_RVT U7070 ( .A1(n12385), .A2(n6759), .Y(n6941) );
  OR2X1_RVT U7071 ( .A1(n12794), .A2(n6547), .Y(n6759) );
  OR2X1_RVT U7072 ( .A1(n7171), .A2(n6708), .Y(n7155) );
  AND2X1_RVT U7073 ( .A1(n6661), .A2(n6933), .Y(n7171) );
  OR2X1_RVT U7074 ( .A1(n6517), .A2(n6606), .Y(n6661) );
  OR2X1_RVT U7075 ( .A1(n7172), .A2(n6597), .Y(n7154) );
  AND2X1_RVT U7076 ( .A1(n6560), .A2(n6562), .Y(n7172) );
  AND4X1_RVT U7077 ( .A1(n7173), .A2(n7174), .A3(n7175), .A4(n7176), .Y(n7146)
         );
  AND4X1_RVT U7078 ( .A1(n7177), .A2(n7178), .A3(n7179), .A4(n7180), .Y(n7176)
         );
  OR2X1_RVT U7079 ( .A1(n7181), .A2(n12388), .Y(n7180) );
  AND2X1_RVT U7080 ( .A1(n6488), .A2(n6780), .Y(n7181) );
  OR2X1_RVT U7081 ( .A1(n6637), .A2(n6668), .Y(n6780) );
  OR2X1_RVT U7082 ( .A1(n12391), .A2(n6520), .Y(n6668) );
  OR2X1_RVT U7083 ( .A1(n12395), .A2(n7182), .Y(n6488) );
  OR2X1_RVT U7084 ( .A1(n12378), .A2(n12384), .Y(n7182) );
  OR2X1_RVT U7085 ( .A1(n7183), .A2(n12402), .Y(n7179) );
  AND2X1_RVT U7086 ( .A1(n6797), .A2(n7184), .Y(n7183) );
  OR2X1_RVT U7087 ( .A1(n12407), .A2(n174), .Y(n7184) );
  OR2X1_RVT U7088 ( .A1(n12405), .A2(n6604), .Y(n6797) );
  OR2X1_RVT U7089 ( .A1(n7185), .A2(n12383), .Y(n7178) );
  AND2X1_RVT U7090 ( .A1(n6815), .A2(n7186), .Y(n7185) );
  OR2X1_RVT U7091 ( .A1(n12408), .A2(n6540), .Y(n7186) );
  OR2X1_RVT U7092 ( .A1(n6482), .A2(n7187), .Y(n6815) );
  OR2X1_RVT U7093 ( .A1(n7188), .A2(n6541), .Y(n7177) );
  AND2X1_RVT U7094 ( .A1(n7189), .A2(n7190), .Y(n7188) );
  OR2X1_RVT U7095 ( .A1(n6597), .A2(n12405), .Y(n7190) );
  AND2X1_RVT U7096 ( .A1(n7191), .A2(n6573), .Y(n7189) );
  OR2X1_RVT U7097 ( .A1(n6559), .A2(n6520), .Y(n6573) );
  OR2X1_RVT U7098 ( .A1(n12380), .A2(n6604), .Y(n7191) );
  OR2X1_RVT U7099 ( .A1(n12802), .A2(n6559), .Y(n6604) );
  OR2X1_RVT U7100 ( .A1(n7192), .A2(n6617), .Y(n7175) );
  AND4X1_RVT U7101 ( .A1(n7193), .A2(n7194), .A3(n6770), .A4(n6680), .Y(n7192)
         );
  OR2X1_RVT U7102 ( .A1(n6743), .A2(n6843), .Y(n6680) );
  OR2X1_RVT U7103 ( .A1(n6575), .A2(n7121), .Y(n6770) );
  OR2X1_RVT U7104 ( .A1(n12386), .A2(n12379), .Y(n7121) );
  OR2X1_RVT U7105 ( .A1(n176), .A2(n6497), .Y(n7194) );
  OR2X1_RVT U7106 ( .A1(n174), .A2(n12405), .Y(n7193) );
  OR2X1_RVT U7107 ( .A1(n7195), .A2(n6553), .Y(n7174) );
  AND2X1_RVT U7108 ( .A1(n7196), .A2(n6574), .Y(n7195) );
  AND2X1_RVT U7109 ( .A1(n7128), .A2(n6824), .Y(n7196) );
  OR2X1_RVT U7110 ( .A1(n7197), .A2(n12799), .Y(n6824) );
  AND2X1_RVT U7111 ( .A1(n6595), .A2(n7198), .Y(n7197) );
  OR2X1_RVT U7112 ( .A1(n12383), .A2(n6482), .Y(n7198) );
  OR2X1_RVT U7113 ( .A1(n6643), .A2(n6781), .Y(n7128) );
  OR2X1_RVT U7114 ( .A1(n6628), .A2(n6517), .Y(n6781) );
  OR2X1_RVT U7115 ( .A1(n7199), .A2(n6621), .Y(n7173) );
  AND2X1_RVT U7116 ( .A1(n7200), .A2(n12391), .Y(n7199) );
  AND2X1_RVT U7117 ( .A1(n7201), .A2(n6802), .Y(n7200) );
  OR2X1_RVT U7118 ( .A1(n6643), .A2(n6743), .Y(n7201) );
  AND4X1_RVT U7119 ( .A1(n7202), .A2(n7203), .A3(n7204), .A4(n7205), .Y(n7145)
         );
  AND2X1_RVT U7120 ( .A1(n7206), .A2(n7207), .Y(n7205) );
  OR2X1_RVT U7121 ( .A1(n12795), .A2(n6723), .Y(n7207) );
  OR2X1_RVT U7122 ( .A1(n12399), .A2(n7208), .Y(n6723) );
  OR2X1_RVT U7123 ( .A1(n6539), .A2(n6628), .Y(n7208) );
  AND2X1_RVT U7124 ( .A1(n7209), .A2(n7210), .Y(n7206) );
  OR2X1_RVT U7125 ( .A1(n6512), .A2(n6523), .Y(n7210) );
  OR2X1_RVT U7126 ( .A1(n6556), .A2(n6751), .Y(n6523) );
  OR2X1_RVT U7127 ( .A1(n12791), .A2(n6517), .Y(n6751) );
  OR2X1_RVT U7128 ( .A1(n6559), .A2(n6636), .Y(n7209) );
  OR2X1_RVT U7129 ( .A1(n6547), .A2(n7211), .Y(n6636) );
  OR2X1_RVT U7130 ( .A1(n6547), .A2(n6727), .Y(n7204) );
  OR2X1_RVT U7131 ( .A1(n176), .A2(n12401), .Y(n6727) );
  OR2X1_RVT U7132 ( .A1(n7212), .A2(n6503), .Y(n7203) );
  AND4X1_RVT U7133 ( .A1(n7213), .A2(n7214), .A3(n7215), .A4(n7216), .Y(n7212)
         );
  OR2X1_RVT U7134 ( .A1(n12789), .A2(n7217), .Y(n7215) );
  OR2X1_RVT U7135 ( .A1(n7218), .A2(n12796), .Y(n7217) );
  AND2X1_RVT U7136 ( .A1(n6554), .A2(n7219), .Y(n7218) );
  OR2X1_RVT U7137 ( .A1(n12394), .A2(n7220), .Y(n7214) );
  OR2X1_RVT U7138 ( .A1(n6860), .A2(n6497), .Y(n7220) );
  OR2X1_RVT U7139 ( .A1(n6480), .A2(n6506), .Y(n7213) );
  OR2X1_RVT U7140 ( .A1(n12793), .A2(n6606), .Y(n6506) );
  OR2X1_RVT U7141 ( .A1(n7079), .A2(n6894), .Y(n7202) );
  OR2X1_RVT U7142 ( .A1(n12410), .A2(n6517), .Y(n6894) );
  AND4X1_RVT U7143 ( .A1(n7222), .A2(n7223), .A3(n7224), .A4(n7225), .Y(n7221)
         );
  AND4X1_RVT U7144 ( .A1(n7226), .A2(n7227), .A3(n7228), .A4(n7229), .Y(n7225)
         );
  AND4X1_RVT U7145 ( .A1(n7230), .A2(n7231), .A3(n7232), .A4(n7233), .Y(n7229)
         );
  OR2X1_RVT U7146 ( .A1(n7067), .A2(n7211), .Y(n7233) );
  OR2X1_RVT U7147 ( .A1(n12792), .A2(n12404), .Y(n7211) );
  OR2X1_RVT U7148 ( .A1(n12378), .A2(n12388), .Y(n7067) );
  OR2X1_RVT U7149 ( .A1(n7234), .A2(n6554), .Y(n7232) );
  AND2X1_RVT U7150 ( .A1(n6500), .A2(n7166), .Y(n7234) );
  OR2X1_RVT U7151 ( .A1(n176), .A2(n7235), .Y(n6500) );
  OR2X1_RVT U7152 ( .A1(n12378), .A2(n12789), .Y(n7235) );
  OR2X1_RVT U7153 ( .A1(n7236), .A2(n6482), .Y(n7231) );
  OR2X1_RVT U7154 ( .A1(n12392), .A2(n6643), .Y(n6482) );
  AND2X1_RVT U7155 ( .A1(n6618), .A2(n7237), .Y(n7236) );
  OR2X1_RVT U7156 ( .A1(n6497), .A2(n6699), .Y(n7237) );
  OR2X1_RVT U7157 ( .A1(n12396), .A2(n12384), .Y(n6497) );
  OR2X1_RVT U7158 ( .A1(n6743), .A2(n7238), .Y(n6618) );
  OR2X1_RVT U7159 ( .A1(n12800), .A2(n12399), .Y(n7238) );
  OR2X1_RVT U7160 ( .A1(n7239), .A2(n6541), .Y(n7230) );
  AND2X1_RVT U7161 ( .A1(n6938), .A2(n7240), .Y(n7239) );
  OR2X1_RVT U7162 ( .A1(n7241), .A2(n12789), .Y(n7240) );
  AND2X1_RVT U7163 ( .A1(n6597), .A2(n6950), .Y(n7241) );
  OR2X1_RVT U7164 ( .A1(n12797), .A2(n6559), .Y(n6950) );
  OR2X1_RVT U7165 ( .A1(n12405), .A2(n7242), .Y(n6938) );
  OR2X1_RVT U7166 ( .A1(n12802), .A2(n12798), .Y(n7242) );
  OR2X1_RVT U7167 ( .A1(n7243), .A2(n12383), .Y(n7228) );
  AND2X1_RVT U7168 ( .A1(n7244), .A2(n7245), .Y(n7243) );
  OR2X1_RVT U7169 ( .A1(n7246), .A2(n6643), .Y(n7245) );
  AND2X1_RVT U7170 ( .A1(n6708), .A2(n7247), .Y(n7246) );
  OR2X1_RVT U7171 ( .A1(n6499), .A2(n6621), .Y(n7244) );
  OR2X1_RVT U7172 ( .A1(n12397), .A2(n6557), .Y(n6621) );
  OR2X1_RVT U7173 ( .A1(n7248), .A2(n12798), .Y(n7227) );
  AND2X1_RVT U7174 ( .A1(n6713), .A2(n6872), .Y(n7248) );
  OR2X1_RVT U7175 ( .A1(n12395), .A2(n7249), .Y(n6872) );
  OR2X1_RVT U7176 ( .A1(n6553), .A2(n12384), .Y(n7249) );
  OR2X1_RVT U7177 ( .A1(n6499), .A2(n7079), .Y(n6713) );
  OR2X1_RVT U7178 ( .A1(n12384), .A2(n12399), .Y(n7079) );
  OR2X1_RVT U7179 ( .A1(n7250), .A2(n12381), .Y(n7226) );
  AND2X1_RVT U7180 ( .A1(n6753), .A2(n7251), .Y(n7250) );
  OR2X1_RVT U7181 ( .A1(n7066), .A2(n6547), .Y(n7251) );
  OR2X1_RVT U7182 ( .A1(n6606), .A2(n7187), .Y(n6753) );
  OR2X1_RVT U7183 ( .A1(n12797), .A2(n176), .Y(n7187) );
  AND2X1_RVT U7184 ( .A1(n12385), .A2(n12800), .Y(n6849) );
  AND4X1_RVT U7185 ( .A1(n7252), .A2(n7253), .A3(n7254), .A4(n7255), .Y(n7224)
         );
  AND4X1_RVT U7186 ( .A1(n7256), .A2(n7257), .A3(n7258), .A4(n7259), .Y(n7255)
         );
  OR2X1_RVT U7187 ( .A1(n7260), .A2(n12390), .Y(n7259) );
  AND2X1_RVT U7188 ( .A1(n6740), .A2(n6811), .Y(n7260) );
  OR2X1_RVT U7189 ( .A1(n6556), .A2(n7166), .Y(n6811) );
  OR2X1_RVT U7190 ( .A1(n12800), .A2(n6553), .Y(n7166) );
  OR2X1_RVT U7191 ( .A1(n12787), .A2(n12380), .Y(n6556) );
  OR2X1_RVT U7192 ( .A1(n12381), .A2(n6843), .Y(n6740) );
  OR2X1_RVT U7193 ( .A1(n12385), .A2(n12399), .Y(n6843) );
  OR2X1_RVT U7194 ( .A1(n7261), .A2(n12796), .Y(n7258) );
  AND2X1_RVT U7195 ( .A1(n6902), .A2(n7262), .Y(n7261) );
  OR2X1_RVT U7196 ( .A1(n6860), .A2(n6570), .Y(n7262) );
  OR2X1_RVT U7197 ( .A1(n6743), .A2(n7263), .Y(n6570) );
  OR2X1_RVT U7198 ( .A1(n12410), .A2(n12386), .Y(n7263) );
  OR2X1_RVT U7199 ( .A1(n12394), .A2(n7264), .Y(n6902) );
  OR2X1_RVT U7200 ( .A1(n6743), .A2(n6539), .Y(n7264) );
  OR2X1_RVT U7201 ( .A1(n7265), .A2(n12802), .Y(n7257) );
  AND2X1_RVT U7202 ( .A1(n6848), .A2(n6777), .Y(n7265) );
  OR2X1_RVT U7203 ( .A1(n6559), .A2(n6595), .Y(n6777) );
  OR2X1_RVT U7204 ( .A1(n12794), .A2(n6743), .Y(n6595) );
  OR2X1_RVT U7205 ( .A1(n7066), .A2(n6575), .Y(n6848) );
  OR2X1_RVT U7206 ( .A1(n12391), .A2(n12799), .Y(n7066) );
  OR2X1_RVT U7207 ( .A1(n7266), .A2(n6617), .Y(n7256) );
  AND2X1_RVT U7208 ( .A1(n7267), .A2(n7268), .Y(n7266) );
  OR2X1_RVT U7209 ( .A1(n6539), .A2(n7065), .Y(n7268) );
  OR2X1_RVT U7210 ( .A1(n12796), .A2(n184), .Y(n7065) );
  AND2X1_RVT U7211 ( .A1(n7269), .A2(n6834), .Y(n7267) );
  OR2X1_RVT U7212 ( .A1(n6547), .A2(n7270), .Y(n6834) );
  OR2X1_RVT U7213 ( .A1(n12407), .A2(n12386), .Y(n7270) );
  OR2X1_RVT U7214 ( .A1(n6603), .A2(n6540), .Y(n7254) );
  OR2X1_RVT U7215 ( .A1(n12789), .A2(n6499), .Y(n6603) );
  OR2X1_RVT U7216 ( .A1(n7271), .A2(n6503), .Y(n7253) );
  AND2X1_RVT U7217 ( .A1(n7272), .A2(n6684), .Y(n7271) );
  AND2X1_RVT U7218 ( .A1(n7273), .A2(n7274), .Y(n6684) );
  OR2X1_RVT U7219 ( .A1(n12395), .A2(n6708), .Y(n7274) );
  OR2X1_RVT U7220 ( .A1(n6606), .A2(n6480), .Y(n7273) );
  OR2X1_RVT U7221 ( .A1(n12380), .A2(n6553), .Y(n6480) );
  AND2X1_RVT U7222 ( .A1(n7275), .A2(n6870), .Y(n7272) );
  OR2X1_RVT U7223 ( .A1(n6637), .A2(n7219), .Y(n6870) );
  OR2X1_RVT U7224 ( .A1(n12791), .A2(n174), .Y(n7219) );
  OR2X1_RVT U7225 ( .A1(n6499), .A2(n6666), .Y(n7275) );
  OR2X1_RVT U7226 ( .A1(n12379), .A2(n7276), .Y(n6666) );
  OR2X1_RVT U7227 ( .A1(n12787), .A2(n12408), .Y(n7276) );
  OR2X1_RVT U7228 ( .A1(n7277), .A2(n12787), .Y(n7252) );
  AND4X1_RVT U7229 ( .A1(n7278), .A2(n7279), .A3(n7280), .A4(n7111), .Y(n7277)
         );
  OR2X1_RVT U7230 ( .A1(n6553), .A2(n6933), .Y(n7111) );
  OR2X1_RVT U7231 ( .A1(n12792), .A2(n12798), .Y(n6933) );
  OR2X1_RVT U7232 ( .A1(n6553), .A2(n7281), .Y(n7280) );
  OR2X1_RVT U7233 ( .A1(n12385), .A2(n12390), .Y(n7281) );
  OR2X1_RVT U7234 ( .A1(n12797), .A2(n6512), .Y(n6553) );
  OR2X1_RVT U7235 ( .A1(n7282), .A2(n6634), .Y(n7279) );
  OR2X1_RVT U7236 ( .A1(n12379), .A2(n6478), .Y(n6634) );
  AND2X1_RVT U7237 ( .A1(n6617), .A2(n7283), .Y(n7282) );
  OR2X1_RVT U7238 ( .A1(n12795), .A2(n6517), .Y(n7283) );
  OR2X1_RVT U7239 ( .A1(n12791), .A2(n12390), .Y(n6617) );
  OR2X1_RVT U7240 ( .A1(n12793), .A2(n7247), .Y(n7278) );
  OR2X1_RVT U7241 ( .A1(n12797), .A2(n6557), .Y(n7247) );
  OR2X1_RVT U7242 ( .A1(n6503), .A2(n174), .Y(n6557) );
  AND4X1_RVT U7243 ( .A1(n7284), .A2(n7285), .A3(n7286), .A4(n7287), .Y(n7223)
         );
  AND4X1_RVT U7244 ( .A1(n7288), .A2(n7289), .A3(n7290), .A4(n7291), .Y(n7287)
         );
  OR2X1_RVT U7245 ( .A1(n6575), .A2(n6702), .Y(n7291) );
  OR2X1_RVT U7246 ( .A1(n12392), .A2(n6597), .Y(n6702) );
  OR2X1_RVT U7247 ( .A1(n12396), .A2(n6743), .Y(n6575) );
  OR2X1_RVT U7248 ( .A1(n6562), .A2(n7137), .Y(n7290) );
  OR2X1_RVT U7249 ( .A1(n12801), .A2(n12379), .Y(n7137) );
  OR2X1_RVT U7250 ( .A1(n6628), .A2(n6554), .Y(n6562) );
  OR2X1_RVT U7251 ( .A1(n6547), .A2(n6574), .Y(n7289) );
  OR2X1_RVT U7252 ( .A1(n12388), .A2(n12401), .Y(n6574) );
  OR2X1_RVT U7253 ( .A1(n12378), .A2(n12788), .Y(n6547) );
  OR2X1_RVT U7254 ( .A1(n184), .A2(n6913), .Y(n7288) );
  OR2X1_RVT U7255 ( .A1(n12386), .A2(n6700), .Y(n6913) );
  OR2X1_RVT U7256 ( .A1(n6517), .A2(n6947), .Y(n7286) );
  OR2X1_RVT U7257 ( .A1(n184), .A2(n7292), .Y(n6947) );
  OR2X1_RVT U7258 ( .A1(n12794), .A2(n12399), .Y(n7292) );
  AND2X1_RVT U7259 ( .A1(n12380), .A2(n12383), .Y(n7076) );
  OR2X1_RVT U7260 ( .A1(n6559), .A2(n6507), .Y(n7285) );
  OR2X1_RVT U7261 ( .A1(n12408), .A2(n7293), .Y(n6507) );
  OR2X1_RVT U7262 ( .A1(n12795), .A2(n12787), .Y(n7293) );
  OR2X1_RVT U7263 ( .A1(n12385), .A2(n6539), .Y(n6559) );
  OR2X1_RVT U7264 ( .A1(n6606), .A2(n7269), .Y(n7284) );
  OR2X1_RVT U7265 ( .A1(n12381), .A2(n6561), .Y(n7269) );
  OR2X1_RVT U7266 ( .A1(n12797), .A2(n12798), .Y(n6561) );
  AND4X1_RVT U7267 ( .A1(n7294), .A2(n6672), .A3(n7295), .A4(n7296), .Y(n7222)
         );
  OR2X1_RVT U7268 ( .A1(n12385), .A2(n7216), .Y(n7296) );
  OR2X1_RVT U7269 ( .A1(n12793), .A2(n6667), .Y(n7216) );
  OR2X1_RVT U7270 ( .A1(n12383), .A2(n6708), .Y(n6667) );
  OR2X1_RVT U7271 ( .A1(n12378), .A2(n6534), .Y(n6708) );
  AND2X1_RVT U7272 ( .A1(n7297), .A2(n7298), .Y(n7295) );
  OR2X1_RVT U7273 ( .A1(n12407), .A2(n7136), .Y(n7298) );
  OR2X1_RVT U7274 ( .A1(n6606), .A2(n6699), .Y(n7136) );
  OR2X1_RVT U7275 ( .A1(n12385), .A2(n12379), .Y(n6699) );
  OR2X1_RVT U7276 ( .A1(n12380), .A2(n6495), .Y(n6534) );
  OR2X1_RVT U7277 ( .A1(n12800), .A2(n6768), .Y(n7297) );
  OR2X1_RVT U7278 ( .A1(n12404), .A2(n6802), .Y(n6768) );
  OR2X1_RVT U7279 ( .A1(n12792), .A2(n12787), .Y(n6802) );
  OR2X1_RVT U7280 ( .A1(n12790), .A2(n12396), .Y(n6478) );
  AND2X1_RVT U7281 ( .A1(n7299), .A2(n7300), .Y(n6672) );
  OR2X1_RVT U7282 ( .A1(n6554), .A2(n6540), .Y(n7300) );
  OR2X1_RVT U7283 ( .A1(n12799), .A2(n6512), .Y(n6540) );
  AND2X1_RVT U7284 ( .A1(n6539), .A2(n6503), .Y(n6592) );
  OR2X1_RVT U7285 ( .A1(n12391), .A2(n6606), .Y(n6554) );
  OR2X1_RVT U7286 ( .A1(n12788), .A2(n6643), .Y(n6606) );
  OR2X1_RVT U7287 ( .A1(n7301), .A2(n6597), .Y(n7299) );
  OR2X1_RVT U7288 ( .A1(n12385), .A2(n174), .Y(n6597) );
  AND2X1_RVT U7289 ( .A1(n12801), .A2(n12378), .Y(n6860) );
  OR2X1_RVT U7290 ( .A1(n12384), .A2(n6700), .Y(n7301) );
  OR2X1_RVT U7291 ( .A1(n12797), .A2(n12401), .Y(n6700) );
  AND2X1_RVT U7292 ( .A1(n7302), .A2(n7303), .Y(n7294) );
  OR2X1_RVT U7293 ( .A1(n6520), .A2(n6853), .Y(n7303) );
  OR2X1_RVT U7294 ( .A1(n12386), .A2(n6560), .Y(n6853) );
  OR2X1_RVT U7295 ( .A1(n12401), .A2(n6637), .Y(n6560) );
  OR2X1_RVT U7296 ( .A1(n12381), .A2(n12384), .Y(n6637) );
  OR2X1_RVT U7297 ( .A1(n12794), .A2(n12792), .Y(n6499) );
  OR2X1_RVT U7298 ( .A1(n12802), .A2(n12796), .Y(n6520) );
  XOR2X1_RVT U7299 ( .A1(key[60]), .A2(state[60]), .Y(n6495) );
  OR2X1_RVT U7300 ( .A1(n6512), .A2(n6641), .Y(n7302) );
  OR2X1_RVT U7301 ( .A1(n6743), .A2(n6934), .Y(n6641) );
  OR2X1_RVT U7302 ( .A1(n12388), .A2(n6541), .Y(n6934) );
  OR2X1_RVT U7303 ( .A1(n12795), .A2(n6643), .Y(n6541) );
  XOR2X1_RVT U7304 ( .A1(key[58]), .A2(state[58]), .Y(n6643) );
  XOR2X1_RVT U7305 ( .A1(key[59]), .A2(state[59]), .Y(n6577) );
  OR2X1_RVT U7306 ( .A1(n12800), .A2(n12386), .Y(n6517) );
  XOR2X1_RVT U7307 ( .A1(key[61]), .A2(state[61]), .Y(n6503) );
  XOR2X1_RVT U7308 ( .A1(key[62]), .A2(state[62]), .Y(n6539) );
  OR2X1_RVT U7309 ( .A1(n12790), .A2(n12384), .Y(n6743) );
  XOR2X1_RVT U7310 ( .A1(key[56]), .A2(state[56]), .Y(n6518) );
  XOR2X1_RVT U7311 ( .A1(key[57]), .A2(state[57]), .Y(n6628) );
  XOR2X1_RVT U7312 ( .A1(key[63]), .A2(state[63]), .Y(n6512) );
  AND4X1_RVT U7313 ( .A1(n7305), .A2(n7306), .A3(n7307), .A4(n7308), .Y(n7304)
         );
  AND4X1_RVT U7314 ( .A1(n7309), .A2(n7310), .A3(n7311), .A4(n7312), .Y(n7308)
         );
  AND4X1_RVT U7315 ( .A1(n7313), .A2(n7314), .A3(n7315), .A4(n7316), .Y(n7312)
         );
  OR2X1_RVT U7316 ( .A1(n12372), .A2(n7318), .Y(n7311) );
  OR2X1_RVT U7317 ( .A1(n7319), .A2(n7320), .Y(n7309) );
  OR2X1_RVT U7318 ( .A1(n12784), .A2(n7321), .Y(n7320) );
  AND4X1_RVT U7319 ( .A1(n7322), .A2(n7323), .A3(n7324), .A4(n7325), .Y(n7307)
         );
  OR2X1_RVT U7320 ( .A1(n7326), .A2(n12782), .Y(n7325) );
  AND2X1_RVT U7321 ( .A1(n7327), .A2(n7328), .Y(n7326) );
  AND2X1_RVT U7322 ( .A1(n7329), .A2(n7330), .Y(n7324) );
  OR2X1_RVT U7323 ( .A1(n7331), .A2(n196), .Y(n7330) );
  AND2X1_RVT U7324 ( .A1(n7332), .A2(n7333), .Y(n7331) );
  OR2X1_RVT U7325 ( .A1(n12363), .A2(n7335), .Y(n7333) );
  OR2X1_RVT U7326 ( .A1(n7321), .A2(n7336), .Y(n7332) );
  OR2X1_RVT U7327 ( .A1(n7337), .A2(n12369), .Y(n7329) );
  AND2X1_RVT U7328 ( .A1(n7339), .A2(n7340), .Y(n7337) );
  OR2X1_RVT U7329 ( .A1(n7341), .A2(n7342), .Y(n7323) );
  AND2X1_RVT U7330 ( .A1(n7343), .A2(n7344), .Y(n7341) );
  OR2X1_RVT U7331 ( .A1(n12364), .A2(n7345), .Y(n7344) );
  AND2X1_RVT U7332 ( .A1(n7346), .A2(n7347), .Y(n7343) );
  AND2X1_RVT U7333 ( .A1(n7348), .A2(n7349), .Y(n7322) );
  OR2X1_RVT U7334 ( .A1(n7350), .A2(n12346), .Y(n7349) );
  AND2X1_RVT U7335 ( .A1(n7352), .A2(n7353), .Y(n7350) );
  OR2X1_RVT U7336 ( .A1(n7354), .A2(n7355), .Y(n7353) );
  OR2X1_RVT U7337 ( .A1(n12355), .A2(n12350), .Y(n7355) );
  OR2X1_RVT U7338 ( .A1(n7358), .A2(n7359), .Y(n7348) );
  AND2X1_RVT U7339 ( .A1(n7360), .A2(n7361), .Y(n7358) );
  AND2X1_RVT U7340 ( .A1(n7362), .A2(n7363), .Y(n7360) );
  AND4X1_RVT U7341 ( .A1(n7364), .A2(n7365), .A3(n7366), .A4(n7367), .Y(n7306)
         );
  AND4X1_RVT U7342 ( .A1(n7368), .A2(n7369), .A3(n7370), .A4(n7371), .Y(n7367)
         );
  OR2X1_RVT U7343 ( .A1(n7372), .A2(n12375), .Y(n7371) );
  AND4X1_RVT U7344 ( .A1(n7374), .A2(n7375), .A3(n7376), .A4(n7377), .Y(n7372)
         );
  OR2X1_RVT U7345 ( .A1(n7378), .A2(n7345), .Y(n7377) );
  OR2X1_RVT U7346 ( .A1(n7379), .A2(n12361), .Y(n7376) );
  OR2X1_RVT U7347 ( .A1(n7381), .A2(n12352), .Y(n7370) );
  AND4X1_RVT U7348 ( .A1(n7382), .A2(n7383), .A3(n7384), .A4(n7385), .Y(n7381)
         );
  OR2X1_RVT U7349 ( .A1(n7386), .A2(n7387), .Y(n7385) );
  OR2X1_RVT U7350 ( .A1(n12369), .A2(n12364), .Y(n7387) );
  AND2X1_RVT U7351 ( .A1(n7388), .A2(n7389), .Y(n7384) );
  OR2X1_RVT U7352 ( .A1(n12786), .A2(n7390), .Y(n7383) );
  OR2X1_RVT U7353 ( .A1(n7391), .A2(n7392), .Y(n7382) );
  AND2X1_RVT U7354 ( .A1(n7393), .A2(n7394), .Y(n7391) );
  OR2X1_RVT U7355 ( .A1(n12369), .A2(n7395), .Y(n7394) );
  OR2X1_RVT U7356 ( .A1(n7328), .A2(n7396), .Y(n7369) );
  OR2X1_RVT U7357 ( .A1(n7395), .A2(n7397), .Y(n7368) );
  OR2X1_RVT U7358 ( .A1(n7398), .A2(n7399), .Y(n7366) );
  OR2X1_RVT U7359 ( .A1(n7400), .A2(n7393), .Y(n7365) );
  OR2X1_RVT U7360 ( .A1(n7401), .A2(n7402), .Y(n7364) );
  AND4X1_RVT U7361 ( .A1(n7403), .A2(n7404), .A3(n7405), .A4(n7406), .Y(n7305)
         );
  AND2X1_RVT U7362 ( .A1(n7407), .A2(n7408), .Y(n7406) );
  OR2X1_RVT U7363 ( .A1(n7392), .A2(n7409), .Y(n7408) );
  AND2X1_RVT U7364 ( .A1(n7410), .A2(n7411), .Y(n7407) );
  OR2X1_RVT U7365 ( .A1(n7412), .A2(n7335), .Y(n7411) );
  OR2X1_RVT U7366 ( .A1(n7336), .A2(n7413), .Y(n7410) );
  OR2X1_RVT U7367 ( .A1(n194), .A2(n7414), .Y(n7405) );
  OR2X1_RVT U7368 ( .A1(n7415), .A2(n12359), .Y(n7404) );
  OR2X1_RVT U7369 ( .A1(n12362), .A2(n7417), .Y(n7403) );
  AND4X1_RVT U7370 ( .A1(n7419), .A2(n7420), .A3(n7421), .A4(n7422), .Y(n7418)
         );
  AND4X1_RVT U7371 ( .A1(n7423), .A2(n7314), .A3(n7424), .A4(n7425), .Y(n7422)
         );
  AND4X1_RVT U7372 ( .A1(n7426), .A2(n7427), .A3(n7428), .A4(n7429), .Y(n7425)
         );
  OR2X1_RVT U7373 ( .A1(n7335), .A2(n7430), .Y(n7429) );
  OR2X1_RVT U7374 ( .A1(n7431), .A2(n12374), .Y(n7430) );
  OR2X1_RVT U7375 ( .A1(n7336), .A2(n7432), .Y(n7428) );
  OR2X1_RVT U7376 ( .A1(n194), .A2(n12358), .Y(n7432) );
  OR2X1_RVT U7377 ( .A1(n7433), .A2(n7379), .Y(n7427) );
  AND2X1_RVT U7378 ( .A1(n7390), .A2(n7434), .Y(n7433) );
  OR2X1_RVT U7379 ( .A1(n7435), .A2(n7436), .Y(n7426) );
  AND2X1_RVT U7380 ( .A1(n7437), .A2(n7438), .Y(n7435) );
  AND2X1_RVT U7381 ( .A1(n7439), .A2(n7440), .Y(n7424) );
  OR2X1_RVT U7382 ( .A1(n7386), .A2(n7441), .Y(n7440) );
  OR2X1_RVT U7383 ( .A1(n7442), .A2(n12784), .Y(n7441) );
  OR2X1_RVT U7384 ( .A1(n7443), .A2(n7444), .Y(n7439) );
  OR2X1_RVT U7385 ( .A1(n7445), .A2(n12363), .Y(n7444) );
  OR2X1_RVT U7386 ( .A1(n7321), .A2(n7446), .Y(n7314) );
  AND4X1_RVT U7387 ( .A1(n7447), .A2(n7448), .A3(n7449), .A4(n7450), .Y(n7421)
         );
  AND4X1_RVT U7388 ( .A1(n7451), .A2(n7452), .A3(n7453), .A4(n7454), .Y(n7450)
         );
  OR2X1_RVT U7389 ( .A1(n7455), .A2(n12377), .Y(n7454) );
  AND2X1_RVT U7390 ( .A1(n7457), .A2(n7458), .Y(n7455) );
  OR2X1_RVT U7391 ( .A1(n12346), .A2(n7336), .Y(n7458) );
  OR2X1_RVT U7392 ( .A1(n7459), .A2(n7338), .Y(n7453) );
  AND2X1_RVT U7393 ( .A1(n7460), .A2(n7461), .Y(n7459) );
  OR2X1_RVT U7394 ( .A1(n7462), .A2(n12783), .Y(n7452) );
  AND2X1_RVT U7395 ( .A1(n7463), .A2(n7464), .Y(n7462) );
  OR2X1_RVT U7396 ( .A1(n7465), .A2(n7414), .Y(n7464) );
  AND2X1_RVT U7397 ( .A1(n12377), .A2(n12361), .Y(n7465) );
  OR2X1_RVT U7398 ( .A1(n7466), .A2(n12347), .Y(n7451) );
  AND2X1_RVT U7399 ( .A1(n7468), .A2(n7469), .Y(n7466) );
  OR2X1_RVT U7400 ( .A1(n7470), .A2(n12353), .Y(n7449) );
  AND2X1_RVT U7401 ( .A1(n7471), .A2(n7472), .Y(n7470) );
  OR2X1_RVT U7402 ( .A1(n12361), .A2(n7473), .Y(n7472) );
  AND2X1_RVT U7403 ( .A1(n7474), .A2(n7475), .Y(n7471) );
  OR2X1_RVT U7404 ( .A1(n7476), .A2(n7477), .Y(n7474) );
  OR2X1_RVT U7405 ( .A1(n7321), .A2(n7392), .Y(n7477) );
  OR2X1_RVT U7406 ( .A1(n7478), .A2(n12780), .Y(n7448) );
  AND2X1_RVT U7407 ( .A1(n7479), .A2(n7480), .Y(n7478) );
  OR2X1_RVT U7408 ( .A1(n7481), .A2(n7482), .Y(n7447) );
  AND2X1_RVT U7409 ( .A1(n7483), .A2(n7484), .Y(n7481) );
  AND2X1_RVT U7410 ( .A1(n7485), .A2(n7486), .Y(n7483) );
  OR2X1_RVT U7411 ( .A1(n196), .A2(n7414), .Y(n7486) );
  OR2X1_RVT U7412 ( .A1(n12371), .A2(n7379), .Y(n7485) );
  AND4X1_RVT U7413 ( .A1(n7487), .A2(n7488), .A3(n7489), .A4(n7490), .Y(n7420)
         );
  AND4X1_RVT U7414 ( .A1(n7491), .A2(n7492), .A3(n7493), .A4(n7494), .Y(n7490)
         );
  OR2X1_RVT U7415 ( .A1(n7414), .A2(n7413), .Y(n7494) );
  OR2X1_RVT U7416 ( .A1(n7345), .A2(n7495), .Y(n7493) );
  OR2X1_RVT U7417 ( .A1(n7378), .A2(n7496), .Y(n7492) );
  OR2X1_RVT U7418 ( .A1(n7321), .A2(n7497), .Y(n7491) );
  AND2X1_RVT U7419 ( .A1(n7498), .A2(n7499), .Y(n7489) );
  OR2X1_RVT U7420 ( .A1(n12372), .A2(n7500), .Y(n7499) );
  OR2X1_RVT U7421 ( .A1(n12351), .A2(n7397), .Y(n7498) );
  OR2X1_RVT U7422 ( .A1(n7501), .A2(n7356), .Y(n7488) );
  AND4X1_RVT U7423 ( .A1(n7502), .A2(n7503), .A3(n7504), .A4(n7505), .Y(n7501)
         );
  OR2X1_RVT U7424 ( .A1(n7506), .A2(n7321), .Y(n7504) );
  OR2X1_RVT U7425 ( .A1(n12772), .A2(n7507), .Y(n7503) );
  OR2X1_RVT U7426 ( .A1(n7508), .A2(n12780), .Y(n7502) );
  AND2X1_RVT U7427 ( .A1(n7399), .A2(n7509), .Y(n7508) );
  OR2X1_RVT U7428 ( .A1(n7401), .A2(n7510), .Y(n7487) );
  AND4X1_RVT U7429 ( .A1(n7511), .A2(n7512), .A3(n7513), .A4(n7514), .Y(n7419)
         );
  AND4X1_RVT U7430 ( .A1(n7515), .A2(n7516), .A3(n7517), .A4(n7518), .Y(n7514)
         );
  OR2X1_RVT U7431 ( .A1(n12776), .A2(n7519), .Y(n7518) );
  OR2X1_RVT U7432 ( .A1(n12777), .A2(n7520), .Y(n7517) );
  OR2X1_RVT U7433 ( .A1(n12774), .A2(n7521), .Y(n7516) );
  OR2X1_RVT U7434 ( .A1(n12345), .A2(n7522), .Y(n7515) );
  OR2X1_RVT U7435 ( .A1(n7523), .A2(n12352), .Y(n7512) );
  AND4X1_RVT U7436 ( .A1(n7525), .A2(n7526), .A3(n7527), .A4(n7528), .Y(n7524)
         );
  AND4X1_RVT U7437 ( .A1(n7529), .A2(n7530), .A3(n7531), .A4(n7532), .Y(n7528)
         );
  AND4X1_RVT U7438 ( .A1(n7533), .A2(n7310), .A3(n7480), .A4(n7534), .Y(n7532)
         );
  OR2X1_RVT U7439 ( .A1(n7535), .A2(n12771), .Y(n7310) );
  AND2X1_RVT U7440 ( .A1(n7536), .A2(n7537), .Y(n7535) );
  OR2X1_RVT U7441 ( .A1(n7354), .A2(n7538), .Y(n7537) );
  OR2X1_RVT U7442 ( .A1(n7539), .A2(n7436), .Y(n7536) );
  OR2X1_RVT U7443 ( .A1(n7540), .A2(n7395), .Y(n7533) );
  AND2X1_RVT U7444 ( .A1(n7541), .A2(n7542), .Y(n7540) );
  OR2X1_RVT U7445 ( .A1(n12776), .A2(n7379), .Y(n7542) );
  OR2X1_RVT U7446 ( .A1(n7543), .A2(n7338), .Y(n7531) );
  AND2X1_RVT U7447 ( .A1(n7544), .A2(n7545), .Y(n7543) );
  OR2X1_RVT U7448 ( .A1(n7546), .A2(n12782), .Y(n7545) );
  AND2X1_RVT U7449 ( .A1(n7386), .A2(n7547), .Y(n7546) );
  OR2X1_RVT U7450 ( .A1(n7548), .A2(n12372), .Y(n7530) );
  AND2X1_RVT U7451 ( .A1(n7549), .A2(n7550), .Y(n7548) );
  OR2X1_RVT U7452 ( .A1(n7379), .A2(n7345), .Y(n7550) );
  OR2X1_RVT U7453 ( .A1(n7551), .A2(n12355), .Y(n7529) );
  AND2X1_RVT U7454 ( .A1(n7463), .A2(n7552), .Y(n7551) );
  OR2X1_RVT U7455 ( .A1(n7392), .A2(n7553), .Y(n7463) );
  AND4X1_RVT U7456 ( .A1(n7554), .A2(n7555), .A3(n7556), .A4(n7557), .Y(n7527)
         );
  OR2X1_RVT U7457 ( .A1(n7558), .A2(n12362), .Y(n7557) );
  AND2X1_RVT U7458 ( .A1(n7559), .A2(n7560), .Y(n7558) );
  OR2X1_RVT U7459 ( .A1(n7436), .A2(n7336), .Y(n7560) );
  AND2X1_RVT U7460 ( .A1(n7561), .A2(n7562), .Y(n7559) );
  OR2X1_RVT U7461 ( .A1(n7476), .A2(n7538), .Y(n7561) );
  AND2X1_RVT U7462 ( .A1(n7563), .A2(n7564), .Y(n7556) );
  OR2X1_RVT U7463 ( .A1(n7565), .A2(n7467), .Y(n7564) );
  AND2X1_RVT U7464 ( .A1(n7566), .A2(n7375), .Y(n7565) );
  OR2X1_RVT U7465 ( .A1(n7321), .A2(n7436), .Y(n7375) );
  OR2X1_RVT U7466 ( .A1(n7567), .A2(n196), .Y(n7563) );
  AND2X1_RVT U7467 ( .A1(n7568), .A2(n7569), .Y(n7567) );
  OR2X1_RVT U7468 ( .A1(n7570), .A2(n12364), .Y(n7569) );
  AND2X1_RVT U7469 ( .A1(n7571), .A2(n7572), .Y(n7570) );
  OR2X1_RVT U7470 ( .A1(n12359), .A2(n7386), .Y(n7572) );
  OR2X1_RVT U7471 ( .A1(n12786), .A2(n12361), .Y(n7571) );
  AND2X1_RVT U7472 ( .A1(n7437), .A2(n7547), .Y(n7568) );
  OR2X1_RVT U7473 ( .A1(n7467), .A2(n7573), .Y(n7437) );
  OR2X1_RVT U7474 ( .A1(n12781), .A2(n12777), .Y(n7573) );
  OR2X1_RVT U7475 ( .A1(n7574), .A2(n7456), .Y(n7555) );
  AND4X1_RVT U7476 ( .A1(n7415), .A2(n7575), .A3(n7576), .A4(n7577), .Y(n7574)
         );
  OR2X1_RVT U7477 ( .A1(n12363), .A2(n7436), .Y(n7577) );
  AND2X1_RVT U7478 ( .A1(n7578), .A2(n7579), .Y(n7576) );
  OR2X1_RVT U7479 ( .A1(n12786), .A2(n12372), .Y(n7575) );
  AND2X1_RVT U7480 ( .A1(n7580), .A2(n7581), .Y(n7415) );
  OR2X1_RVT U7481 ( .A1(n7582), .A2(n194), .Y(n7581) );
  OR2X1_RVT U7482 ( .A1(n7379), .A2(n12771), .Y(n7580) );
  AND2X1_RVT U7483 ( .A1(n7583), .A2(n7584), .Y(n7554) );
  OR2X1_RVT U7484 ( .A1(n7585), .A2(n12773), .Y(n7584) );
  AND2X1_RVT U7485 ( .A1(n7586), .A2(n7587), .Y(n7585) );
  OR2X1_RVT U7486 ( .A1(n7588), .A2(n12366), .Y(n7587) );
  AND2X1_RVT U7487 ( .A1(n7589), .A2(n7590), .Y(n7588) );
  AND2X1_RVT U7488 ( .A1(n7591), .A2(n7592), .Y(n7586) );
  OR2X1_RVT U7489 ( .A1(n7593), .A2(n12375), .Y(n7583) );
  AND4X1_RVT U7490 ( .A1(n7594), .A2(n7595), .A3(n7596), .A4(n7597), .Y(n7593)
         );
  OR2X1_RVT U7491 ( .A1(n12785), .A2(n7598), .Y(n7596) );
  OR2X1_RVT U7492 ( .A1(n194), .A2(n7393), .Y(n7595) );
  OR2X1_RVT U7493 ( .A1(n7482), .A2(n7436), .Y(n7594) );
  AND4X1_RVT U7494 ( .A1(n7599), .A2(n7600), .A3(n7601), .A4(n7602), .Y(n7526)
         );
  AND2X1_RVT U7495 ( .A1(n7603), .A2(n7446), .Y(n7602) );
  OR2X1_RVT U7496 ( .A1(n12350), .A2(n7412), .Y(n7446) );
  AND2X1_RVT U7497 ( .A1(n7604), .A2(n7605), .Y(n7603) );
  OR2X1_RVT U7498 ( .A1(n7606), .A2(n7361), .Y(n7605) );
  OR2X1_RVT U7499 ( .A1(n7413), .A2(n7473), .Y(n7604) );
  OR2X1_RVT U7500 ( .A1(n194), .A2(n7607), .Y(n7601) );
  OR2X1_RVT U7501 ( .A1(n12784), .A2(n7608), .Y(n7600) );
  OR2X1_RVT U7502 ( .A1(n7482), .A2(n7609), .Y(n7599) );
  AND4X1_RVT U7503 ( .A1(n7610), .A2(n7611), .A3(n7612), .A4(n7613), .Y(n7525)
         );
  AND2X1_RVT U7504 ( .A1(n7614), .A2(n7615), .Y(n7613) );
  OR2X1_RVT U7505 ( .A1(n12345), .A2(n7616), .Y(n7615) );
  AND2X1_RVT U7506 ( .A1(n7617), .A2(n7618), .Y(n7614) );
  OR2X1_RVT U7507 ( .A1(n7378), .A2(n7388), .Y(n7618) );
  OR2X1_RVT U7508 ( .A1(n12366), .A2(n7438), .Y(n7388) );
  OR2X1_RVT U7509 ( .A1(n12352), .A2(n7619), .Y(n7617) );
  OR2X1_RVT U7510 ( .A1(n7359), .A2(n7352), .Y(n7612) );
  OR2X1_RVT U7511 ( .A1(n7445), .A2(n7620), .Y(n7352) );
  OR2X1_RVT U7512 ( .A1(n12780), .A2(n7621), .Y(n7611) );
  OR2X1_RVT U7513 ( .A1(n12364), .A2(n7479), .Y(n7610) );
  OR2X1_RVT U7514 ( .A1(n12771), .A2(n7541), .Y(n7479) );
  AND4X1_RVT U7515 ( .A1(n7623), .A2(n7624), .A3(n7625), .A4(n7626), .Y(n7622)
         );
  AND4X1_RVT U7516 ( .A1(n7627), .A2(n7628), .A3(n7629), .A4(n7630), .Y(n7626)
         );
  OR2X1_RVT U7517 ( .A1(n204), .A2(n7631), .Y(n7630) );
  OR2X1_RVT U7518 ( .A1(n7632), .A2(n12377), .Y(n7631) );
  AND2X1_RVT U7519 ( .A1(n12366), .A2(n7398), .Y(n7632) );
  AND2X1_RVT U7520 ( .A1(n7313), .A2(n7633), .Y(n7629) );
  OR2X1_RVT U7521 ( .A1(n12355), .A2(n7634), .Y(n7313) );
  OR2X1_RVT U7522 ( .A1(n204), .A2(n7392), .Y(n7634) );
  OR2X1_RVT U7523 ( .A1(n7635), .A2(n7321), .Y(n7628) );
  AND2X1_RVT U7524 ( .A1(n7636), .A2(n7637), .Y(n7635) );
  AND2X1_RVT U7525 ( .A1(n7638), .A2(n7639), .Y(n7627) );
  OR2X1_RVT U7526 ( .A1(n7640), .A2(n7641), .Y(n7639) );
  AND2X1_RVT U7527 ( .A1(n7642), .A2(n7402), .Y(n7640) );
  OR2X1_RVT U7528 ( .A1(n7643), .A2(n7393), .Y(n7638) );
  AND2X1_RVT U7529 ( .A1(n7578), .A2(n7412), .Y(n7643) );
  OR2X1_RVT U7530 ( .A1(n12353), .A2(n7644), .Y(n7578) );
  OR2X1_RVT U7531 ( .A1(n12786), .A2(n12363), .Y(n7644) );
  AND4X1_RVT U7532 ( .A1(n7645), .A2(n7646), .A3(n7647), .A4(n7648), .Y(n7625)
         );
  OR2X1_RVT U7533 ( .A1(n7649), .A2(n12776), .Y(n7648) );
  AND2X1_RVT U7534 ( .A1(n7461), .A2(n7650), .Y(n7649) );
  OR2X1_RVT U7535 ( .A1(n12784), .A2(n7506), .Y(n7461) );
  AND2X1_RVT U7536 ( .A1(n7651), .A2(n7652), .Y(n7647) );
  OR2X1_RVT U7537 ( .A1(n7653), .A2(n12774), .Y(n7652) );
  AND2X1_RVT U7538 ( .A1(n7654), .A2(n7655), .Y(n7653) );
  OR2X1_RVT U7539 ( .A1(n7356), .A2(n7598), .Y(n7655) );
  OR2X1_RVT U7540 ( .A1(n7656), .A2(n12772), .Y(n7651) );
  AND2X1_RVT U7541 ( .A1(n7657), .A2(n7658), .Y(n7656) );
  OR2X1_RVT U7542 ( .A1(n7659), .A2(n12366), .Y(n7646) );
  AND2X1_RVT U7543 ( .A1(n7660), .A2(n7661), .Y(n7659) );
  AND2X1_RVT U7544 ( .A1(n7662), .A2(n7663), .Y(n7660) );
  AND2X1_RVT U7545 ( .A1(n7664), .A2(n7665), .Y(n7645) );
  OR2X1_RVT U7546 ( .A1(n7666), .A2(n7582), .Y(n7665) );
  AND2X1_RVT U7547 ( .A1(n7667), .A2(n7413), .Y(n7666) );
  AND2X1_RVT U7548 ( .A1(n7668), .A2(n7669), .Y(n7667) );
  OR2X1_RVT U7549 ( .A1(n7670), .A2(n12369), .Y(n7664) );
  AND2X1_RVT U7550 ( .A1(n7671), .A2(n7672), .Y(n7670) );
  OR2X1_RVT U7551 ( .A1(n12783), .A2(n12371), .Y(n7672) );
  AND2X1_RVT U7552 ( .A1(n7402), .A2(n7673), .Y(n7671) );
  AND4X1_RVT U7553 ( .A1(n7674), .A2(n7675), .A3(n7676), .A4(n7677), .Y(n7624)
         );
  AND2X1_RVT U7554 ( .A1(n7678), .A2(n7679), .Y(n7677) );
  OR2X1_RVT U7555 ( .A1(n7395), .A2(n7469), .Y(n7679) );
  OR2X1_RVT U7556 ( .A1(n12778), .A2(n7402), .Y(n7469) );
  AND2X1_RVT U7557 ( .A1(n7680), .A2(n7681), .Y(n7678) );
  OR2X1_RVT U7558 ( .A1(n7547), .A2(n7361), .Y(n7681) );
  OR2X1_RVT U7559 ( .A1(n12785), .A2(n12362), .Y(n7361) );
  OR2X1_RVT U7560 ( .A1(n7445), .A2(n7495), .Y(n7680) );
  OR2X1_RVT U7561 ( .A1(n12773), .A2(n7682), .Y(n7495) );
  OR2X1_RVT U7562 ( .A1(n7683), .A2(n12345), .Y(n7676) );
  AND4X1_RVT U7563 ( .A1(n7684), .A2(n7685), .A3(n7686), .A4(n7687), .Y(n7683)
         );
  OR2X1_RVT U7564 ( .A1(n7620), .A2(n7393), .Y(n7686) );
  OR2X1_RVT U7565 ( .A1(n7688), .A2(n7390), .Y(n7685) );
  OR2X1_RVT U7566 ( .A1(n12782), .A2(n7345), .Y(n7684) );
  OR2X1_RVT U7567 ( .A1(n7689), .A2(n12346), .Y(n7675) );
  AND2X1_RVT U7568 ( .A1(n7690), .A2(n7691), .Y(n7689) );
  OR2X1_RVT U7569 ( .A1(n7620), .A2(n7345), .Y(n7691) );
  AND2X1_RVT U7570 ( .A1(n7692), .A2(n7621), .Y(n7690) );
  OR2X1_RVT U7571 ( .A1(n7393), .A2(n7693), .Y(n7621) );
  OR2X1_RVT U7572 ( .A1(n12773), .A2(n12785), .Y(n7693) );
  OR2X1_RVT U7573 ( .A1(n7694), .A2(n12353), .Y(n7674) );
  AND4X1_RVT U7574 ( .A1(n7695), .A2(n7608), .A3(n7417), .A4(n7389), .Y(n7694)
         );
  OR2X1_RVT U7575 ( .A1(n7414), .A2(n7696), .Y(n7389) );
  OR2X1_RVT U7576 ( .A1(n12775), .A2(n7351), .Y(n7696) );
  OR2X1_RVT U7577 ( .A1(n7476), .A2(n7510), .Y(n7417) );
  OR2X1_RVT U7578 ( .A1(n7395), .A2(n7697), .Y(n7608) );
  OR2X1_RVT U7579 ( .A1(n12377), .A2(n12346), .Y(n7697) );
  OR2X1_RVT U7580 ( .A1(n7354), .A2(n7698), .Y(n7695) );
  OR2X1_RVT U7581 ( .A1(n7699), .A2(n12351), .Y(n7698) );
  AND4X1_RVT U7582 ( .A1(n7700), .A2(n7701), .A3(n7702), .A4(n7703), .Y(n7623)
         );
  AND2X1_RVT U7583 ( .A1(n7704), .A2(n7705), .Y(n7703) );
  AND2X1_RVT U7584 ( .A1(n7706), .A2(n7707), .Y(n7704) );
  OR2X1_RVT U7585 ( .A1(n7386), .A2(n7661), .Y(n7707) );
  OR2X1_RVT U7586 ( .A1(n7398), .A2(n7708), .Y(n7661) );
  OR2X1_RVT U7587 ( .A1(n12774), .A2(n12776), .Y(n7708) );
  OR2X1_RVT U7588 ( .A1(n12781), .A2(n7709), .Y(n7706) );
  OR2X1_RVT U7589 ( .A1(n12362), .A2(n7710), .Y(n7702) );
  OR2X1_RVT U7590 ( .A1(n12784), .A2(n7711), .Y(n7701) );
  OR2X1_RVT U7591 ( .A1(n7398), .A2(n7712), .Y(n7700) );
  AND4X1_RVT U7592 ( .A1(n7714), .A2(n7715), .A3(n7716), .A4(n7717), .Y(n7713)
         );
  AND4X1_RVT U7593 ( .A1(n7718), .A2(n7719), .A3(n7720), .A4(n7721), .Y(n7717)
         );
  AND4X1_RVT U7594 ( .A1(n7722), .A2(n7723), .A3(n7315), .A4(n7724), .Y(n7721)
         );
  OR2X1_RVT U7595 ( .A1(n7456), .A2(n7725), .Y(n7315) );
  OR2X1_RVT U7596 ( .A1(n7547), .A2(n196), .Y(n7725) );
  OR2X1_RVT U7597 ( .A1(n7319), .A2(n7726), .Y(n7723) );
  OR2X1_RVT U7598 ( .A1(n12779), .A2(n12782), .Y(n7726) );
  OR2X1_RVT U7599 ( .A1(n7582), .A2(n7727), .Y(n7722) );
  OR2X1_RVT U7600 ( .A1(n7728), .A2(n7356), .Y(n7727) );
  AND2X1_RVT U7601 ( .A1(n12366), .A2(n7456), .Y(n7728) );
  OR2X1_RVT U7602 ( .A1(n7729), .A2(n12372), .Y(n7720) );
  AND2X1_RVT U7603 ( .A1(n7597), .A2(n7669), .Y(n7729) );
  OR2X1_RVT U7604 ( .A1(n196), .A2(n7730), .Y(n7669) );
  OR2X1_RVT U7605 ( .A1(n12345), .A2(n12778), .Y(n7730) );
  OR2X1_RVT U7606 ( .A1(n7386), .A2(n7731), .Y(n7597) );
  OR2X1_RVT U7607 ( .A1(n12776), .A2(n7378), .Y(n7731) );
  OR2X1_RVT U7608 ( .A1(n7732), .A2(n7336), .Y(n7719) );
  AND2X1_RVT U7609 ( .A1(n7733), .A2(n7541), .Y(n7732) );
  OR2X1_RVT U7610 ( .A1(n7442), .A2(n7436), .Y(n7718) );
  AND4X1_RVT U7611 ( .A1(n7734), .A2(n7735), .A3(n7736), .A4(n7737), .Y(n7716)
         );
  AND2X1_RVT U7612 ( .A1(n7738), .A2(n7739), .Y(n7737) );
  OR2X1_RVT U7613 ( .A1(n7740), .A2(n12366), .Y(n7739) );
  AND2X1_RVT U7614 ( .A1(n7741), .A2(n7409), .Y(n7740) );
  AND2X1_RVT U7615 ( .A1(n7742), .A2(n7743), .Y(n7738) );
  OR2X1_RVT U7616 ( .A1(n7744), .A2(n7392), .Y(n7743) );
  AND2X1_RVT U7617 ( .A1(n7363), .A2(n7335), .Y(n7744) );
  OR2X1_RVT U7618 ( .A1(n12784), .A2(n7434), .Y(n7363) );
  OR2X1_RVT U7619 ( .A1(n7745), .A2(n7445), .Y(n7742) );
  AND2X1_RVT U7620 ( .A1(n7637), .A2(n7746), .Y(n7745) );
  OR2X1_RVT U7621 ( .A1(n12785), .A2(n7473), .Y(n7637) );
  OR2X1_RVT U7622 ( .A1(n7747), .A2(n12776), .Y(n7736) );
  AND2X1_RVT U7623 ( .A1(n7340), .A2(n7748), .Y(n7747) );
  OR2X1_RVT U7624 ( .A1(n7476), .A2(n7400), .Y(n7748) );
  OR2X1_RVT U7625 ( .A1(n7379), .A2(n7582), .Y(n7340) );
  OR2X1_RVT U7626 ( .A1(n7749), .A2(n194), .Y(n7735) );
  AND2X1_RVT U7627 ( .A1(n7390), .A2(n7750), .Y(n7749) );
  OR2X1_RVT U7628 ( .A1(n7751), .A2(n12350), .Y(n7750) );
  AND2X1_RVT U7629 ( .A1(n7752), .A2(n7753), .Y(n7751) );
  OR2X1_RVT U7630 ( .A1(n12777), .A2(n7373), .Y(n7753) );
  OR2X1_RVT U7631 ( .A1(n12377), .A2(n7476), .Y(n7390) );
  OR2X1_RVT U7632 ( .A1(n7754), .A2(n7460), .Y(n7734) );
  AND2X1_RVT U7633 ( .A1(n7393), .A2(n7438), .Y(n7754) );
  OR2X1_RVT U7634 ( .A1(n12773), .A2(n7321), .Y(n7438) );
  AND4X1_RVT U7635 ( .A1(n7755), .A2(n7756), .A3(n7757), .A4(n7758), .Y(n7715)
         );
  AND4X1_RVT U7636 ( .A1(n7759), .A2(n7760), .A3(n7761), .A4(n7762), .Y(n7758)
         );
  OR2X1_RVT U7637 ( .A1(n7763), .A2(n12784), .Y(n7762) );
  AND2X1_RVT U7638 ( .A1(n7496), .A2(n7764), .Y(n7763) );
  OR2X1_RVT U7639 ( .A1(n12374), .A2(n7345), .Y(n7764) );
  OR2X1_RVT U7640 ( .A1(n7765), .A2(n7338), .Y(n7761) );
  AND2X1_RVT U7641 ( .A1(n7766), .A2(n7767), .Y(n7765) );
  OR2X1_RVT U7642 ( .A1(n7768), .A2(n7373), .Y(n7767) );
  AND2X1_RVT U7643 ( .A1(n7398), .A2(n7386), .Y(n7768) );
  AND2X1_RVT U7644 ( .A1(n7400), .A2(n7642), .Y(n7766) );
  OR2X1_RVT U7645 ( .A1(n12375), .A2(n7538), .Y(n7642) );
  OR2X1_RVT U7646 ( .A1(n7769), .A2(n12364), .Y(n7760) );
  AND2X1_RVT U7647 ( .A1(n7770), .A2(n7771), .Y(n7769) );
  OR2X1_RVT U7648 ( .A1(n7386), .A2(n7772), .Y(n7771) );
  AND2X1_RVT U7649 ( .A1(n7468), .A2(n7662), .Y(n7770) );
  OR2X1_RVT U7650 ( .A1(n7378), .A2(n7553), .Y(n7662) );
  OR2X1_RVT U7651 ( .A1(n7351), .A2(n7773), .Y(n7468) );
  OR2X1_RVT U7652 ( .A1(n7774), .A2(n7321), .Y(n7759) );
  AND4X1_RVT U7653 ( .A1(n7775), .A2(n7776), .A3(n7777), .A4(n7710), .Y(n7774)
         );
  OR2X1_RVT U7654 ( .A1(n7414), .A2(n7778), .Y(n7710) );
  OR2X1_RVT U7655 ( .A1(n12345), .A2(n7378), .Y(n7778) );
  OR2X1_RVT U7656 ( .A1(n12781), .A2(n7620), .Y(n7776) );
  OR2X1_RVT U7657 ( .A1(n7379), .A2(n7476), .Y(n7775) );
  OR2X1_RVT U7658 ( .A1(n7547), .A2(n7589), .Y(n7757) );
  OR2X1_RVT U7659 ( .A1(n7779), .A2(n12348), .Y(n7756) );
  AND4X1_RVT U7660 ( .A1(n7780), .A2(n7781), .A3(n7423), .A4(n7521), .Y(n7779)
         );
  OR2X1_RVT U7661 ( .A1(n7345), .A2(n7510), .Y(n7521) );
  OR2X1_RVT U7662 ( .A1(n12781), .A2(n194), .Y(n7510) );
  OR2X1_RVT U7663 ( .A1(n7338), .A2(n7402), .Y(n7423) );
  OR2X1_RVT U7664 ( .A1(n12773), .A2(n7773), .Y(n7755) );
  AND4X1_RVT U7665 ( .A1(n7782), .A2(n7783), .A3(n7784), .A4(n7785), .Y(n7714)
         );
  OR2X1_RVT U7666 ( .A1(n12353), .A2(n7786), .Y(n7785) );
  AND2X1_RVT U7667 ( .A1(n7787), .A2(n7788), .Y(n7784) );
  OR2X1_RVT U7668 ( .A1(n12374), .A2(n7541), .Y(n7788) );
  OR2X1_RVT U7669 ( .A1(n7328), .A2(n7402), .Y(n7787) );
  OR2X1_RVT U7670 ( .A1(n196), .A2(n7359), .Y(n7402) );
  OR2X1_RVT U7671 ( .A1(n12377), .A2(n7520), .Y(n7783) );
  OR2X1_RVT U7672 ( .A1(n7395), .A2(n7789), .Y(n7520) );
  AND2X1_RVT U7673 ( .A1(n7790), .A2(n7791), .Y(n7782) );
  OR2X1_RVT U7674 ( .A1(n12346), .A2(n7792), .Y(n7791) );
  OR2X1_RVT U7675 ( .A1(n7398), .A2(n7347), .Y(n7790) );
  OR2X1_RVT U7676 ( .A1(n7321), .A2(n7606), .Y(n7347) );
  AND4X1_RVT U7677 ( .A1(n7794), .A2(n7795), .A3(n7796), .A4(n7797), .Y(n7793)
         );
  AND4X1_RVT U7678 ( .A1(n7798), .A2(n7799), .A3(n7800), .A4(n7801), .Y(n7797)
         );
  AND4X1_RVT U7679 ( .A1(n7534), .A2(n7724), .A3(n7802), .A4(n7803), .Y(n7801)
         );
  OR2X1_RVT U7680 ( .A1(n7804), .A2(n7805), .Y(n7724) );
  OR2X1_RVT U7681 ( .A1(n7319), .A2(n7589), .Y(n7534) );
  OR2X1_RVT U7682 ( .A1(n12782), .A2(n12362), .Y(n7589) );
  AND4X1_RVT U7683 ( .A1(n7792), .A2(n7658), .A3(n7781), .A4(n7316), .Y(n7800)
         );
  OR2X1_RVT U7684 ( .A1(n7806), .A2(n7506), .Y(n7316) );
  OR2X1_RVT U7685 ( .A1(n7321), .A2(n7807), .Y(n7781) );
  OR2X1_RVT U7686 ( .A1(n7354), .A2(n194), .Y(n7658) );
  OR2X1_RVT U7687 ( .A1(n7345), .A2(n7808), .Y(n7792) );
  OR2X1_RVT U7688 ( .A1(n12352), .A2(n12372), .Y(n7808) );
  AND4X1_RVT U7689 ( .A1(n7809), .A2(n7810), .A3(n7811), .A4(n7812), .Y(n7799)
         );
  OR2X1_RVT U7690 ( .A1(n7598), .A2(n7813), .Y(n7812) );
  OR2X1_RVT U7691 ( .A1(n12372), .A2(n7378), .Y(n7813) );
  OR2X1_RVT U7692 ( .A1(n7507), .A2(n7814), .Y(n7811) );
  OR2X1_RVT U7693 ( .A1(n12783), .A2(n7395), .Y(n7814) );
  OR2X1_RVT U7694 ( .A1(n7733), .A2(n7815), .Y(n7810) );
  OR2X1_RVT U7695 ( .A1(n7816), .A2(n7392), .Y(n7815) );
  OR2X1_RVT U7696 ( .A1(n12369), .A2(n7817), .Y(n7809) );
  OR2X1_RVT U7697 ( .A1(n7818), .A2(n12352), .Y(n7817) );
  AND2X1_RVT U7698 ( .A1(n7606), .A2(n7819), .Y(n7818) );
  AND2X1_RVT U7699 ( .A1(n7820), .A2(n7821), .Y(n7798) );
  OR2X1_RVT U7700 ( .A1(n7822), .A2(n7373), .Y(n7821) );
  AND2X1_RVT U7701 ( .A1(n7823), .A2(n7824), .Y(n7822) );
  OR2X1_RVT U7702 ( .A1(n12351), .A2(n7566), .Y(n7824) );
  OR2X1_RVT U7703 ( .A1(n12355), .A2(n7641), .Y(n7823) );
  AND2X1_RVT U7704 ( .A1(n7825), .A2(n7826), .Y(n7820) );
  OR2X1_RVT U7705 ( .A1(n7827), .A2(n7412), .Y(n7826) );
  AND2X1_RVT U7706 ( .A1(n7828), .A2(n7829), .Y(n7827) );
  OR2X1_RVT U7707 ( .A1(n12358), .A2(n204), .Y(n7829) );
  NAND2X1_RVT U7708 ( .A1(n7395), .A2(n12775), .Y(n7828) );
  OR2X1_RVT U7709 ( .A1(n7830), .A2(n196), .Y(n7825) );
  AND2X1_RVT U7710 ( .A1(n7619), .A2(n7496), .Y(n7830) );
  OR2X1_RVT U7711 ( .A1(n7345), .A2(n7831), .Y(n7496) );
  OR2X1_RVT U7712 ( .A1(n12786), .A2(n12347), .Y(n7831) );
  AND4X1_RVT U7713 ( .A1(n7513), .A2(n7832), .A3(n7705), .A4(n7833), .Y(n7796)
         );
  AND4X1_RVT U7714 ( .A1(n7834), .A2(n7835), .A3(n7836), .A4(n7837), .Y(n7833)
         );
  OR2X1_RVT U7715 ( .A1(n7476), .A2(n7397), .Y(n7837) );
  OR2X1_RVT U7716 ( .A1(n7414), .A2(n7443), .Y(n7836) );
  OR2X1_RVT U7717 ( .A1(n12774), .A2(n7668), .Y(n7835) );
  OR2X1_RVT U7718 ( .A1(n7392), .A2(n7374), .Y(n7668) );
  OR2X1_RVT U7719 ( .A1(n12782), .A2(n7456), .Y(n7374) );
  OR2X1_RVT U7720 ( .A1(n12361), .A2(n7497), .Y(n7834) );
  OR2X1_RVT U7721 ( .A1(n7378), .A2(n7606), .Y(n7497) );
  OR2X1_RVT U7722 ( .A1(n12345), .A2(n7582), .Y(n7606) );
  AND2X1_RVT U7723 ( .A1(n7838), .A2(n7839), .Y(n7705) );
  OR2X1_RVT U7724 ( .A1(n7840), .A2(n7445), .Y(n7839) );
  OR2X1_RVT U7725 ( .A1(n12371), .A2(n196), .Y(n7840) );
  OR2X1_RVT U7726 ( .A1(n7841), .A2(n7328), .Y(n7838) );
  OR2X1_RVT U7727 ( .A1(n12773), .A2(n7445), .Y(n7328) );
  OR2X1_RVT U7728 ( .A1(n7342), .A2(n7392), .Y(n7841) );
  OR2X1_RVT U7729 ( .A1(n12353), .A2(n7711), .Y(n7832) );
  AND2X1_RVT U7730 ( .A1(n7842), .A2(n7843), .Y(n7513) );
  OR2X1_RVT U7731 ( .A1(n7396), .A2(n7434), .Y(n7843) );
  OR2X1_RVT U7732 ( .A1(n7844), .A2(n7845), .Y(n7842) );
  AND4X1_RVT U7733 ( .A1(n7846), .A2(n7847), .A3(n7848), .A4(n7849), .Y(n7795)
         );
  OR2X1_RVT U7734 ( .A1(n7850), .A2(n7582), .Y(n7849) );
  AND2X1_RVT U7735 ( .A1(n7851), .A2(n7591), .Y(n7850) );
  OR2X1_RVT U7736 ( .A1(n12359), .A2(n7807), .Y(n7591) );
  OR2X1_RVT U7737 ( .A1(n7852), .A2(n12779), .Y(n7848) );
  AND2X1_RVT U7738 ( .A1(n7519), .A2(n7484), .Y(n7852) );
  OR2X1_RVT U7739 ( .A1(n12773), .A2(n7460), .Y(n7484) );
  OR2X1_RVT U7740 ( .A1(n7853), .A2(n7539), .Y(n7847) );
  AND2X1_RVT U7741 ( .A1(n7854), .A2(n7855), .Y(n7853) );
  OR2X1_RVT U7742 ( .A1(n12348), .A2(n7398), .Y(n7855) );
  AND2X1_RVT U7743 ( .A1(n7856), .A2(n7436), .Y(n7854) );
  OR2X1_RVT U7744 ( .A1(n194), .A2(n7395), .Y(n7856) );
  OR2X1_RVT U7745 ( .A1(n7857), .A2(n7336), .Y(n7846) );
  AND2X1_RVT U7746 ( .A1(n7858), .A2(n7859), .Y(n7857) );
  NAND2X1_RVT U7747 ( .A1(n7321), .A2(n7699), .Y(n7859) );
  AND2X1_RVT U7748 ( .A1(n7860), .A2(n7549), .Y(n7858) );
  OR2X1_RVT U7749 ( .A1(n7482), .A2(n7807), .Y(n7549) );
  OR2X1_RVT U7750 ( .A1(n12368), .A2(n7861), .Y(n7860) );
  AND4X1_RVT U7751 ( .A1(n7862), .A2(n7863), .A3(n7864), .A4(n7865), .Y(n7794)
         );
  OR2X1_RVT U7752 ( .A1(n7866), .A2(n7359), .Y(n7865) );
  AND2X1_RVT U7753 ( .A1(n7867), .A2(n7500), .Y(n7866) );
  AND2X1_RVT U7754 ( .A1(n7868), .A2(n7522), .Y(n7867) );
  OR2X1_RVT U7755 ( .A1(n196), .A2(n7845), .Y(n7522) );
  OR2X1_RVT U7756 ( .A1(n12347), .A2(n7456), .Y(n7845) );
  OR2X1_RVT U7757 ( .A1(n7869), .A2(n12364), .Y(n7864) );
  AND2X1_RVT U7758 ( .A1(n7870), .A2(n7871), .Y(n7869) );
  OR2X1_RVT U7759 ( .A1(n7872), .A2(n12771), .Y(n7871) );
  AND2X1_RVT U7760 ( .A1(n7873), .A2(n7874), .Y(n7872) );
  OR2X1_RVT U7761 ( .A1(n12346), .A2(n7733), .Y(n7874) );
  OR2X1_RVT U7762 ( .A1(n12778), .A2(n7379), .Y(n7873) );
  AND2X1_RVT U7763 ( .A1(n7875), .A2(n7876), .Y(n7870) );
  OR2X1_RVT U7764 ( .A1(n7345), .A2(n7877), .Y(n7875) );
  OR2X1_RVT U7765 ( .A1(n7878), .A2(n7379), .Y(n7863) );
  AND4X1_RVT U7766 ( .A1(n7879), .A2(n7880), .A3(n7881), .A4(n7345), .Y(n7878)
         );
  OR2X1_RVT U7767 ( .A1(n12779), .A2(n7395), .Y(n7881) );
  OR2X1_RVT U7768 ( .A1(n12358), .A2(n7414), .Y(n7880) );
  OR2X1_RVT U7769 ( .A1(n7467), .A2(n7445), .Y(n7879) );
  OR2X1_RVT U7770 ( .A1(n7882), .A2(n7321), .Y(n7862) );
  AND4X1_RVT U7771 ( .A1(n7746), .A2(n7883), .A3(n7544), .A4(n7460), .Y(n7882)
         );
  OR2X1_RVT U7772 ( .A1(n7414), .A2(n7877), .Y(n7544) );
  OR2X1_RVT U7773 ( .A1(n7582), .A2(n7789), .Y(n7883) );
  OR2X1_RVT U7774 ( .A1(n12352), .A2(n7547), .Y(n7746) );
  AND4X1_RVT U7775 ( .A1(n7885), .A2(n7886), .A3(n7887), .A4(n7888), .Y(n7884)
         );
  AND4X1_RVT U7776 ( .A1(n7397), .A2(n7633), .A3(n7889), .A4(n7890), .Y(n7888)
         );
  AND4X1_RVT U7777 ( .A1(n7712), .A2(n7657), .A3(n7802), .A4(n7803), .Y(n7890)
         );
  OR2X1_RVT U7778 ( .A1(n7805), .A2(n7318), .Y(n7803) );
  OR2X1_RVT U7779 ( .A1(n12777), .A2(n7436), .Y(n7318) );
  OR2X1_RVT U7780 ( .A1(n7335), .A2(n7844), .Y(n7802) );
  OR2X1_RVT U7781 ( .A1(n12782), .A2(n12366), .Y(n7844) );
  OR2X1_RVT U7782 ( .A1(n12771), .A2(n7456), .Y(n7335) );
  OR2X1_RVT U7783 ( .A1(n12783), .A2(n7354), .Y(n7657) );
  OR2X1_RVT U7784 ( .A1(n12375), .A2(n12359), .Y(n7354) );
  OR2X1_RVT U7785 ( .A1(n7476), .A2(n7891), .Y(n7712) );
  OR2X1_RVT U7786 ( .A1(n12366), .A2(n7380), .Y(n7891) );
  OR2X1_RVT U7787 ( .A1(n7378), .A2(n7892), .Y(n7889) );
  OR2X1_RVT U7788 ( .A1(n7506), .A2(n12357), .Y(n7892) );
  OR2X1_RVT U7789 ( .A1(n7445), .A2(n7893), .Y(n7633) );
  OR2X1_RVT U7790 ( .A1(n7379), .A2(n12364), .Y(n7893) );
  OR2X1_RVT U7791 ( .A1(n12775), .A2(n7804), .Y(n7397) );
  OR2X1_RVT U7792 ( .A1(n12359), .A2(n7396), .Y(n7804) );
  AND4X1_RVT U7793 ( .A1(n7894), .A2(n7895), .A3(n7896), .A4(n7897), .Y(n7887)
         );
  AND4X1_RVT U7794 ( .A1(n7898), .A2(n7899), .A3(n7900), .A4(n7901), .Y(n7897)
         );
  OR2X1_RVT U7795 ( .A1(n7412), .A2(n7902), .Y(n7901) );
  OR2X1_RVT U7796 ( .A1(n12348), .A2(n7482), .Y(n7902) );
  OR2X1_RVT U7797 ( .A1(n7395), .A2(n7903), .Y(n7900) );
  OR2X1_RVT U7798 ( .A1(n7904), .A2(n7359), .Y(n7903) );
  AND2X1_RVT U7799 ( .A1(n7338), .A2(n7398), .Y(n7904) );
  OR2X1_RVT U7800 ( .A1(n7905), .A2(n7906), .Y(n7899) );
  AND2X1_RVT U7801 ( .A1(n7553), .A2(n7509), .Y(n7905) );
  OR2X1_RVT U7802 ( .A1(n12776), .A2(n204), .Y(n7509) );
  OR2X1_RVT U7803 ( .A1(n12772), .A2(n12369), .Y(n7553) );
  OR2X1_RVT U7804 ( .A1(n7907), .A2(n7393), .Y(n7898) );
  AND2X1_RVT U7805 ( .A1(n7789), .A2(n7908), .Y(n7907) );
  OR2X1_RVT U7806 ( .A1(n12774), .A2(n196), .Y(n7908) );
  OR2X1_RVT U7807 ( .A1(n7909), .A2(n12371), .Y(n7896) );
  AND2X1_RVT U7808 ( .A1(n7780), .A2(n7910), .Y(n7909) );
  OR2X1_RVT U7809 ( .A1(n7386), .A2(n7733), .Y(n7910) );
  OR2X1_RVT U7810 ( .A1(n12352), .A2(n7598), .Y(n7780) );
  OR2X1_RVT U7811 ( .A1(n12778), .A2(n7386), .Y(n7598) );
  OR2X1_RVT U7812 ( .A1(n7911), .A2(n7547), .Y(n7895) );
  AND2X1_RVT U7813 ( .A1(n7500), .A2(n7772), .Y(n7911) );
  OR2X1_RVT U7814 ( .A1(n7356), .A2(n7445), .Y(n7500) );
  OR2X1_RVT U7815 ( .A1(n7912), .A2(n7436), .Y(n7894) );
  AND2X1_RVT U7816 ( .A1(n7399), .A2(n7401), .Y(n7912) );
  AND4X1_RVT U7817 ( .A1(n7913), .A2(n7914), .A3(n7915), .A4(n7916), .Y(n7886)
         );
  AND4X1_RVT U7818 ( .A1(n7917), .A2(n7918), .A3(n7919), .A4(n7920), .Y(n7916)
         );
  OR2X1_RVT U7819 ( .A1(n7921), .A2(n12355), .Y(n7920) );
  AND2X1_RVT U7820 ( .A1(n7327), .A2(n7619), .Y(n7921) );
  OR2X1_RVT U7821 ( .A1(n7476), .A2(n7507), .Y(n7619) );
  OR2X1_RVT U7822 ( .A1(n12358), .A2(n7359), .Y(n7507) );
  OR2X1_RVT U7823 ( .A1(n12362), .A2(n7922), .Y(n7327) );
  OR2X1_RVT U7824 ( .A1(n12345), .A2(n12351), .Y(n7922) );
  OR2X1_RVT U7825 ( .A1(n7923), .A2(n12369), .Y(n7919) );
  AND2X1_RVT U7826 ( .A1(n7636), .A2(n7924), .Y(n7923) );
  OR2X1_RVT U7827 ( .A1(n12374), .A2(n194), .Y(n7924) );
  OR2X1_RVT U7828 ( .A1(n12372), .A2(n7443), .Y(n7636) );
  OR2X1_RVT U7829 ( .A1(n7925), .A2(n12350), .Y(n7918) );
  AND2X1_RVT U7830 ( .A1(n7654), .A2(n7926), .Y(n7925) );
  OR2X1_RVT U7831 ( .A1(n12375), .A2(n7379), .Y(n7926) );
  OR2X1_RVT U7832 ( .A1(n7321), .A2(n7927), .Y(n7654) );
  OR2X1_RVT U7833 ( .A1(n7928), .A2(n7380), .Y(n7917) );
  AND2X1_RVT U7834 ( .A1(n7929), .A2(n7930), .Y(n7928) );
  OR2X1_RVT U7835 ( .A1(n7436), .A2(n12372), .Y(n7930) );
  AND2X1_RVT U7836 ( .A1(n7931), .A2(n7412), .Y(n7929) );
  OR2X1_RVT U7837 ( .A1(n7398), .A2(n7359), .Y(n7412) );
  OR2X1_RVT U7838 ( .A1(n12347), .A2(n7443), .Y(n7931) );
  OR2X1_RVT U7839 ( .A1(n12786), .A2(n7398), .Y(n7443) );
  OR2X1_RVT U7840 ( .A1(n7932), .A2(n7456), .Y(n7915) );
  AND4X1_RVT U7841 ( .A1(n7933), .A2(n7934), .A3(n7609), .A4(n7519), .Y(n7932)
         );
  OR2X1_RVT U7842 ( .A1(n7582), .A2(n7682), .Y(n7519) );
  OR2X1_RVT U7843 ( .A1(n7414), .A2(n7861), .Y(n7609) );
  OR2X1_RVT U7844 ( .A1(n12353), .A2(n12346), .Y(n7861) );
  OR2X1_RVT U7845 ( .A1(n196), .A2(n7336), .Y(n7934) );
  OR2X1_RVT U7846 ( .A1(n194), .A2(n12372), .Y(n7933) );
  OR2X1_RVT U7847 ( .A1(n7935), .A2(n7392), .Y(n7914) );
  AND2X1_RVT U7848 ( .A1(n7936), .A2(n7413), .Y(n7935) );
  AND2X1_RVT U7849 ( .A1(n7868), .A2(n7663), .Y(n7936) );
  OR2X1_RVT U7850 ( .A1(n7937), .A2(n12783), .Y(n7663) );
  AND2X1_RVT U7851 ( .A1(n7434), .A2(n7938), .Y(n7937) );
  OR2X1_RVT U7852 ( .A1(n12350), .A2(n7321), .Y(n7938) );
  OR2X1_RVT U7853 ( .A1(n7482), .A2(n7620), .Y(n7868) );
  OR2X1_RVT U7854 ( .A1(n7467), .A2(n7356), .Y(n7620) );
  OR2X1_RVT U7855 ( .A1(n7939), .A2(n7460), .Y(n7913) );
  AND2X1_RVT U7856 ( .A1(n7940), .A2(n12358), .Y(n7939) );
  AND2X1_RVT U7857 ( .A1(n7941), .A2(n7641), .Y(n7940) );
  OR2X1_RVT U7858 ( .A1(n7482), .A2(n7582), .Y(n7941) );
  AND4X1_RVT U7859 ( .A1(n7942), .A2(n7943), .A3(n7944), .A4(n7945), .Y(n7885)
         );
  AND2X1_RVT U7860 ( .A1(n7946), .A2(n7947), .Y(n7945) );
  OR2X1_RVT U7861 ( .A1(n12779), .A2(n7562), .Y(n7947) );
  OR2X1_RVT U7862 ( .A1(n12366), .A2(n7948), .Y(n7562) );
  OR2X1_RVT U7863 ( .A1(n7378), .A2(n7467), .Y(n7948) );
  AND2X1_RVT U7864 ( .A1(n7949), .A2(n7950), .Y(n7946) );
  OR2X1_RVT U7865 ( .A1(n7351), .A2(n7362), .Y(n7950) );
  OR2X1_RVT U7866 ( .A1(n7395), .A2(n7590), .Y(n7362) );
  OR2X1_RVT U7867 ( .A1(n12775), .A2(n7356), .Y(n7590) );
  OR2X1_RVT U7868 ( .A1(n7398), .A2(n7475), .Y(n7949) );
  OR2X1_RVT U7869 ( .A1(n7386), .A2(n7951), .Y(n7475) );
  OR2X1_RVT U7870 ( .A1(n7386), .A2(n7566), .Y(n7944) );
  OR2X1_RVT U7871 ( .A1(n196), .A2(n12368), .Y(n7566) );
  OR2X1_RVT U7872 ( .A1(n7952), .A2(n7342), .Y(n7943) );
  AND4X1_RVT U7873 ( .A1(n7953), .A2(n7954), .A3(n7955), .A4(n7956), .Y(n7952)
         );
  OR2X1_RVT U7874 ( .A1(n12773), .A2(n7957), .Y(n7955) );
  OR2X1_RVT U7875 ( .A1(n7958), .A2(n12780), .Y(n7957) );
  AND2X1_RVT U7876 ( .A1(n7393), .A2(n7959), .Y(n7958) );
  OR2X1_RVT U7877 ( .A1(n12361), .A2(n7960), .Y(n7954) );
  OR2X1_RVT U7878 ( .A1(n7699), .A2(n7336), .Y(n7960) );
  OR2X1_RVT U7879 ( .A1(n7319), .A2(n7345), .Y(n7953) );
  OR2X1_RVT U7880 ( .A1(n12777), .A2(n7445), .Y(n7345) );
  OR2X1_RVT U7881 ( .A1(n7819), .A2(n7733), .Y(n7942) );
  OR2X1_RVT U7882 ( .A1(n12377), .A2(n7356), .Y(n7733) );
  AND4X1_RVT U7883 ( .A1(n7962), .A2(n7963), .A3(n7964), .A4(n7965), .Y(n7961)
         );
  AND4X1_RVT U7884 ( .A1(n7966), .A2(n7967), .A3(n7968), .A4(n7969), .Y(n7965)
         );
  AND4X1_RVT U7885 ( .A1(n7970), .A2(n7971), .A3(n7972), .A4(n7973), .Y(n7969)
         );
  OR2X1_RVT U7886 ( .A1(n7807), .A2(n7951), .Y(n7973) );
  OR2X1_RVT U7887 ( .A1(n12776), .A2(n12371), .Y(n7951) );
  OR2X1_RVT U7888 ( .A1(n12345), .A2(n12355), .Y(n7807) );
  OR2X1_RVT U7889 ( .A1(n7974), .A2(n7393), .Y(n7972) );
  AND2X1_RVT U7890 ( .A1(n7339), .A2(n7906), .Y(n7974) );
  OR2X1_RVT U7891 ( .A1(n196), .A2(n7975), .Y(n7339) );
  OR2X1_RVT U7892 ( .A1(n12345), .A2(n12773), .Y(n7975) );
  OR2X1_RVT U7893 ( .A1(n7976), .A2(n7321), .Y(n7971) );
  OR2X1_RVT U7894 ( .A1(n12359), .A2(n7482), .Y(n7321) );
  AND2X1_RVT U7895 ( .A1(n7457), .A2(n7977), .Y(n7976) );
  OR2X1_RVT U7896 ( .A1(n7336), .A2(n7538), .Y(n7977) );
  OR2X1_RVT U7897 ( .A1(n12363), .A2(n12351), .Y(n7336) );
  OR2X1_RVT U7898 ( .A1(n7582), .A2(n7978), .Y(n7457) );
  OR2X1_RVT U7899 ( .A1(n12784), .A2(n12366), .Y(n7978) );
  OR2X1_RVT U7900 ( .A1(n7979), .A2(n7380), .Y(n7970) );
  AND2X1_RVT U7901 ( .A1(n7777), .A2(n7980), .Y(n7979) );
  OR2X1_RVT U7902 ( .A1(n7981), .A2(n12773), .Y(n7980) );
  AND2X1_RVT U7903 ( .A1(n7436), .A2(n7789), .Y(n7981) );
  OR2X1_RVT U7904 ( .A1(n12781), .A2(n7398), .Y(n7789) );
  OR2X1_RVT U7905 ( .A1(n12372), .A2(n7982), .Y(n7777) );
  OR2X1_RVT U7906 ( .A1(n12786), .A2(n12782), .Y(n7982) );
  OR2X1_RVT U7907 ( .A1(n7983), .A2(n12350), .Y(n7968) );
  AND2X1_RVT U7908 ( .A1(n7984), .A2(n7985), .Y(n7983) );
  OR2X1_RVT U7909 ( .A1(n7986), .A2(n7482), .Y(n7985) );
  AND2X1_RVT U7910 ( .A1(n7547), .A2(n7987), .Y(n7986) );
  OR2X1_RVT U7911 ( .A1(n7338), .A2(n7460), .Y(n7984) );
  OR2X1_RVT U7912 ( .A1(n12364), .A2(n7396), .Y(n7460) );
  OR2X1_RVT U7913 ( .A1(n7988), .A2(n12782), .Y(n7967) );
  AND2X1_RVT U7914 ( .A1(n7552), .A2(n7711), .Y(n7988) );
  OR2X1_RVT U7915 ( .A1(n12362), .A2(n7989), .Y(n7711) );
  OR2X1_RVT U7916 ( .A1(n7392), .A2(n12351), .Y(n7989) );
  OR2X1_RVT U7917 ( .A1(n7338), .A2(n7819), .Y(n7552) );
  OR2X1_RVT U7918 ( .A1(n12351), .A2(n12366), .Y(n7819) );
  OR2X1_RVT U7919 ( .A1(n7990), .A2(n12348), .Y(n7966) );
  AND2X1_RVT U7920 ( .A1(n7592), .A2(n7991), .Y(n7990) );
  OR2X1_RVT U7921 ( .A1(n7806), .A2(n7386), .Y(n7991) );
  OR2X1_RVT U7922 ( .A1(n7445), .A2(n7927), .Y(n7592) );
  OR2X1_RVT U7923 ( .A1(n12781), .A2(n196), .Y(n7927) );
  AND2X1_RVT U7924 ( .A1(n12352), .A2(n12784), .Y(n7688) );
  AND4X1_RVT U7925 ( .A1(n7992), .A2(n7993), .A3(n7994), .A4(n7995), .Y(n7964)
         );
  AND4X1_RVT U7926 ( .A1(n7996), .A2(n7997), .A3(n7998), .A4(n7999), .Y(n7995)
         );
  OR2X1_RVT U7927 ( .A1(n8000), .A2(n12357), .Y(n7999) );
  AND2X1_RVT U7928 ( .A1(n7579), .A2(n7650), .Y(n8000) );
  OR2X1_RVT U7929 ( .A1(n7395), .A2(n7906), .Y(n7650) );
  OR2X1_RVT U7930 ( .A1(n12784), .A2(n7392), .Y(n7906) );
  OR2X1_RVT U7931 ( .A1(n12771), .A2(n12347), .Y(n7395) );
  OR2X1_RVT U7932 ( .A1(n12348), .A2(n7682), .Y(n7579) );
  OR2X1_RVT U7933 ( .A1(n12352), .A2(n12366), .Y(n7682) );
  OR2X1_RVT U7934 ( .A1(n8001), .A2(n12780), .Y(n7998) );
  AND2X1_RVT U7935 ( .A1(n7741), .A2(n8002), .Y(n8001) );
  OR2X1_RVT U7936 ( .A1(n7699), .A2(n7409), .Y(n8002) );
  OR2X1_RVT U7937 ( .A1(n7582), .A2(n8003), .Y(n7409) );
  OR2X1_RVT U7938 ( .A1(n12377), .A2(n12353), .Y(n8003) );
  OR2X1_RVT U7939 ( .A1(n12361), .A2(n8004), .Y(n7741) );
  OR2X1_RVT U7940 ( .A1(n7582), .A2(n7378), .Y(n8004) );
  OR2X1_RVT U7941 ( .A1(n8005), .A2(n12786), .Y(n7997) );
  AND2X1_RVT U7942 ( .A1(n7687), .A2(n7616), .Y(n8005) );
  OR2X1_RVT U7943 ( .A1(n7398), .A2(n7434), .Y(n7616) );
  OR2X1_RVT U7944 ( .A1(n12778), .A2(n7582), .Y(n7434) );
  OR2X1_RVT U7945 ( .A1(n7806), .A2(n7414), .Y(n7687) );
  OR2X1_RVT U7946 ( .A1(n12358), .A2(n12783), .Y(n7806) );
  OR2X1_RVT U7947 ( .A1(n8006), .A2(n7456), .Y(n7996) );
  AND2X1_RVT U7948 ( .A1(n8007), .A2(n8008), .Y(n8006) );
  OR2X1_RVT U7949 ( .A1(n7378), .A2(n7805), .Y(n8008) );
  OR2X1_RVT U7950 ( .A1(n12780), .A2(n204), .Y(n7805) );
  AND2X1_RVT U7951 ( .A1(n8009), .A2(n7673), .Y(n8007) );
  OR2X1_RVT U7952 ( .A1(n7386), .A2(n8010), .Y(n7673) );
  OR2X1_RVT U7953 ( .A1(n12374), .A2(n12353), .Y(n8010) );
  OR2X1_RVT U7954 ( .A1(n7442), .A2(n7379), .Y(n7994) );
  OR2X1_RVT U7955 ( .A1(n12773), .A2(n7338), .Y(n7442) );
  OR2X1_RVT U7956 ( .A1(n8011), .A2(n7342), .Y(n7993) );
  AND2X1_RVT U7957 ( .A1(n8012), .A2(n7523), .Y(n8011) );
  AND2X1_RVT U7958 ( .A1(n8013), .A2(n8014), .Y(n7523) );
  OR2X1_RVT U7959 ( .A1(n12362), .A2(n7547), .Y(n8014) );
  OR2X1_RVT U7960 ( .A1(n7445), .A2(n7319), .Y(n8013) );
  OR2X1_RVT U7961 ( .A1(n12347), .A2(n7392), .Y(n7319) );
  AND2X1_RVT U7962 ( .A1(n8015), .A2(n7709), .Y(n8012) );
  OR2X1_RVT U7963 ( .A1(n7476), .A2(n7959), .Y(n7709) );
  OR2X1_RVT U7964 ( .A1(n12775), .A2(n194), .Y(n7959) );
  OR2X1_RVT U7965 ( .A1(n7338), .A2(n7505), .Y(n8015) );
  OR2X1_RVT U7966 ( .A1(n12346), .A2(n8016), .Y(n7505) );
  OR2X1_RVT U7967 ( .A1(n12771), .A2(n12375), .Y(n8016) );
  OR2X1_RVT U7968 ( .A1(n8017), .A2(n12771), .Y(n7992) );
  AND4X1_RVT U7969 ( .A1(n8018), .A2(n8019), .A3(n8020), .A4(n7851), .Y(n8017)
         );
  OR2X1_RVT U7970 ( .A1(n7392), .A2(n7772), .Y(n7851) );
  OR2X1_RVT U7971 ( .A1(n12776), .A2(n12782), .Y(n7772) );
  OR2X1_RVT U7972 ( .A1(n7392), .A2(n8021), .Y(n8020) );
  OR2X1_RVT U7973 ( .A1(n12352), .A2(n12357), .Y(n8021) );
  OR2X1_RVT U7974 ( .A1(n12781), .A2(n7351), .Y(n7392) );
  OR2X1_RVT U7975 ( .A1(n8022), .A2(n7473), .Y(n8019) );
  OR2X1_RVT U7976 ( .A1(n12346), .A2(n7317), .Y(n7473) );
  AND2X1_RVT U7977 ( .A1(n7456), .A2(n8023), .Y(n8022) );
  OR2X1_RVT U7978 ( .A1(n12779), .A2(n7356), .Y(n8023) );
  OR2X1_RVT U7979 ( .A1(n12775), .A2(n12357), .Y(n7456) );
  OR2X1_RVT U7980 ( .A1(n12777), .A2(n7987), .Y(n8018) );
  OR2X1_RVT U7981 ( .A1(n12781), .A2(n7396), .Y(n7987) );
  OR2X1_RVT U7982 ( .A1(n7342), .A2(n194), .Y(n7396) );
  AND4X1_RVT U7983 ( .A1(n8024), .A2(n8025), .A3(n8026), .A4(n8027), .Y(n7963)
         );
  AND4X1_RVT U7984 ( .A1(n8028), .A2(n8029), .A3(n8030), .A4(n8031), .Y(n8027)
         );
  OR2X1_RVT U7985 ( .A1(n7414), .A2(n7541), .Y(n8031) );
  OR2X1_RVT U7986 ( .A1(n12359), .A2(n7436), .Y(n7541) );
  OR2X1_RVT U7987 ( .A1(n12363), .A2(n7582), .Y(n7414) );
  OR2X1_RVT U7988 ( .A1(n7401), .A2(n7877), .Y(n8030) );
  OR2X1_RVT U7989 ( .A1(n12785), .A2(n12346), .Y(n7877) );
  OR2X1_RVT U7990 ( .A1(n7467), .A2(n7393), .Y(n7401) );
  OR2X1_RVT U7991 ( .A1(n7386), .A2(n7413), .Y(n8029) );
  OR2X1_RVT U7992 ( .A1(n12355), .A2(n12368), .Y(n7413) );
  OR2X1_RVT U7993 ( .A1(n12345), .A2(n12772), .Y(n7386) );
  OR2X1_RVT U7994 ( .A1(n204), .A2(n7752), .Y(n8028) );
  OR2X1_RVT U7995 ( .A1(n12353), .A2(n7539), .Y(n7752) );
  OR2X1_RVT U7996 ( .A1(n7356), .A2(n7786), .Y(n8026) );
  OR2X1_RVT U7997 ( .A1(n204), .A2(n8032), .Y(n7786) );
  OR2X1_RVT U7998 ( .A1(n12778), .A2(n12366), .Y(n8032) );
  AND2X1_RVT U7999 ( .A1(n12347), .A2(n12350), .Y(n7816) );
  OR2X1_RVT U8000 ( .A1(n7398), .A2(n7346), .Y(n8025) );
  OR2X1_RVT U8001 ( .A1(n12375), .A2(n8033), .Y(n7346) );
  OR2X1_RVT U8002 ( .A1(n12779), .A2(n12771), .Y(n8033) );
  OR2X1_RVT U8003 ( .A1(n12352), .A2(n7378), .Y(n7398) );
  OR2X1_RVT U8004 ( .A1(n7445), .A2(n8009), .Y(n8024) );
  OR2X1_RVT U8005 ( .A1(n12348), .A2(n7400), .Y(n8009) );
  OR2X1_RVT U8006 ( .A1(n12781), .A2(n12782), .Y(n7400) );
  AND4X1_RVT U8007 ( .A1(n8034), .A2(n7511), .A3(n8035), .A4(n8036), .Y(n7962)
         );
  OR2X1_RVT U8008 ( .A1(n12352), .A2(n7956), .Y(n8036) );
  OR2X1_RVT U8009 ( .A1(n12777), .A2(n7506), .Y(n7956) );
  OR2X1_RVT U8010 ( .A1(n12350), .A2(n7547), .Y(n7506) );
  OR2X1_RVT U8011 ( .A1(n12345), .A2(n7373), .Y(n7547) );
  AND2X1_RVT U8012 ( .A1(n8037), .A2(n8038), .Y(n8035) );
  OR2X1_RVT U8013 ( .A1(n12374), .A2(n7876), .Y(n8038) );
  OR2X1_RVT U8014 ( .A1(n7445), .A2(n7538), .Y(n7876) );
  OR2X1_RVT U8015 ( .A1(n12352), .A2(n12346), .Y(n7538) );
  OR2X1_RVT U8016 ( .A1(n12347), .A2(n7334), .Y(n7373) );
  OR2X1_RVT U8017 ( .A1(n12784), .A2(n7607), .Y(n8037) );
  OR2X1_RVT U8018 ( .A1(n12371), .A2(n7641), .Y(n7607) );
  OR2X1_RVT U8019 ( .A1(n12776), .A2(n12771), .Y(n7641) );
  OR2X1_RVT U8020 ( .A1(n12774), .A2(n12363), .Y(n7317) );
  AND2X1_RVT U8021 ( .A1(n8039), .A2(n8040), .Y(n7511) );
  OR2X1_RVT U8022 ( .A1(n7393), .A2(n7379), .Y(n8040) );
  OR2X1_RVT U8023 ( .A1(n12783), .A2(n7351), .Y(n7379) );
  AND2X1_RVT U8024 ( .A1(n7378), .A2(n7342), .Y(n7431) );
  OR2X1_RVT U8025 ( .A1(n12358), .A2(n7445), .Y(n7393) );
  OR2X1_RVT U8026 ( .A1(n12772), .A2(n7482), .Y(n7445) );
  OR2X1_RVT U8027 ( .A1(n8041), .A2(n7436), .Y(n8039) );
  OR2X1_RVT U8028 ( .A1(n12352), .A2(n194), .Y(n7436) );
  AND2X1_RVT U8029 ( .A1(n12785), .A2(n12345), .Y(n7699) );
  OR2X1_RVT U8030 ( .A1(n12351), .A2(n7539), .Y(n8041) );
  OR2X1_RVT U8031 ( .A1(n12781), .A2(n12368), .Y(n7539) );
  AND2X1_RVT U8032 ( .A1(n8042), .A2(n8043), .Y(n8034) );
  OR2X1_RVT U8033 ( .A1(n7359), .A2(n7692), .Y(n8043) );
  OR2X1_RVT U8034 ( .A1(n12353), .A2(n7399), .Y(n7692) );
  OR2X1_RVT U8035 ( .A1(n12368), .A2(n7476), .Y(n7399) );
  OR2X1_RVT U8036 ( .A1(n12348), .A2(n12351), .Y(n7476) );
  OR2X1_RVT U8037 ( .A1(n12778), .A2(n12776), .Y(n7338) );
  OR2X1_RVT U8038 ( .A1(n12786), .A2(n12780), .Y(n7359) );
  XOR2X1_RVT U8039 ( .A1(key[52]), .A2(state[52]), .Y(n7334) );
  OR2X1_RVT U8040 ( .A1(n7351), .A2(n7480), .Y(n8042) );
  OR2X1_RVT U8041 ( .A1(n7582), .A2(n7773), .Y(n7480) );
  OR2X1_RVT U8042 ( .A1(n12355), .A2(n7380), .Y(n7773) );
  OR2X1_RVT U8043 ( .A1(n12779), .A2(n7482), .Y(n7380) );
  XOR2X1_RVT U8044 ( .A1(key[50]), .A2(state[50]), .Y(n7482) );
  XOR2X1_RVT U8045 ( .A1(key[51]), .A2(state[51]), .Y(n7416) );
  OR2X1_RVT U8046 ( .A1(n12784), .A2(n12353), .Y(n7356) );
  XOR2X1_RVT U8047 ( .A1(key[53]), .A2(state[53]), .Y(n7342) );
  XOR2X1_RVT U8048 ( .A1(key[54]), .A2(state[54]), .Y(n7378) );
  OR2X1_RVT U8049 ( .A1(n12774), .A2(n12351), .Y(n7582) );
  XOR2X1_RVT U8050 ( .A1(key[48]), .A2(state[48]), .Y(n7357) );
  XOR2X1_RVT U8051 ( .A1(key[49]), .A2(state[49]), .Y(n7467) );
  XOR2X1_RVT U8052 ( .A1(key[55]), .A2(state[55]), .Y(n7351) );
  AND4X1_RVT U8053 ( .A1(n8045), .A2(n8046), .A3(n8047), .A4(n8048), .Y(n8044)
         );
  AND4X1_RVT U8054 ( .A1(n8049), .A2(n8050), .A3(n8051), .A4(n8052), .Y(n8048)
         );
  AND4X1_RVT U8055 ( .A1(n8053), .A2(n1298), .A3(n6124), .A4(n8054), .Y(n8052)
         );
  OR2X1_RVT U8056 ( .A1(n12198), .A2(n7048), .Y(n6124) );
  OR2X1_RVT U8057 ( .A1(n79), .A2(n8055), .Y(n7048) );
  OR2X1_RVT U8058 ( .A1(n8056), .A2(n6132), .Y(n1298) );
  OR2X1_RVT U8059 ( .A1(n76), .A2(n8057), .Y(n8051) );
  OR2X1_RVT U8060 ( .A1(n8058), .A2(n1307), .Y(n8057) );
  AND2X1_RVT U8061 ( .A1(n8059), .A2(n8060), .Y(n8058) );
  OR2X1_RVT U8062 ( .A1(n12190), .A2(n12206), .Y(n8060) );
  OR2X1_RVT U8063 ( .A1(n12877), .A2(n12869), .Y(n8059) );
  OR2X1_RVT U8064 ( .A1(n8061), .A2(n8062), .Y(n8050) );
  OR2X1_RVT U8065 ( .A1(n12150), .A2(n8063), .Y(n8062) );
  OR2X1_RVT U8066 ( .A1(n1348), .A2(n8064), .Y(n8049) );
  OR2X1_RVT U8067 ( .A1(n8065), .A2(n85), .Y(n8064) );
  AND4X1_RVT U8068 ( .A1(n8066), .A2(n8067), .A3(n8068), .A4(n8069), .Y(n8047)
         );
  AND4X1_RVT U8069 ( .A1(n8070), .A2(n8071), .A3(n8072), .A4(n8073), .Y(n8069)
         );
  OR2X1_RVT U8070 ( .A1(n8074), .A2(n1391), .Y(n8073) );
  AND2X1_RVT U8071 ( .A1(n6184), .A2(n7000), .Y(n8074) );
  OR2X1_RVT U8072 ( .A1(n8075), .A2(n12199), .Y(n8072) );
  AND2X1_RVT U8073 ( .A1(n6200), .A2(n6149), .Y(n8075) );
  OR2X1_RVT U8074 ( .A1(n8076), .A2(n12208), .Y(n8071) );
  AND2X1_RVT U8075 ( .A1(n1366), .A2(n8077), .Y(n8076) );
  OR2X1_RVT U8076 ( .A1(n1325), .A2(n8078), .Y(n1366) );
  OR2X1_RVT U8077 ( .A1(n12874), .A2(n85), .Y(n8078) );
  OR2X1_RVT U8078 ( .A1(n8079), .A2(n1356), .Y(n8070) );
  AND2X1_RVT U8079 ( .A1(n6209), .A2(n8080), .Y(n8079) );
  OR2X1_RVT U8080 ( .A1(n6145), .A2(n1306), .Y(n6209) );
  OR2X1_RVT U8081 ( .A1(n8081), .A2(n73), .Y(n8068) );
  AND2X1_RVT U8082 ( .A1(n8082), .A2(n8083), .Y(n8081) );
  OR2X1_RVT U8083 ( .A1(n8084), .A2(n69), .Y(n8067) );
  AND2X1_RVT U8084 ( .A1(n1359), .A2(n1331), .Y(n8084) );
  OR2X1_RVT U8085 ( .A1(n8085), .A2(n12186), .Y(n8066) );
  AND2X1_RVT U8086 ( .A1(n1367), .A2(n8086), .Y(n8085) );
  OR2X1_RVT U8087 ( .A1(n1332), .A2(n8087), .Y(n8086) );
  OR2X1_RVT U8088 ( .A1(n12873), .A2(n12201), .Y(n8087) );
  OR2X1_RVT U8089 ( .A1(n12198), .A2(n8088), .Y(n1367) );
  AND4X1_RVT U8090 ( .A1(n8089), .A2(n8090), .A3(n8091), .A4(n8092), .Y(n8046)
         );
  AND4X1_RVT U8091 ( .A1(n8093), .A2(n8094), .A3(n8095), .A4(n8096), .Y(n8092)
         );
  OR2X1_RVT U8092 ( .A1(n8097), .A2(n12926), .Y(n8096) );
  AND2X1_RVT U8093 ( .A1(n8098), .A2(n8099), .Y(n8097) );
  OR2X1_RVT U8094 ( .A1(n8100), .A2(n1390), .Y(n8099) );
  AND2X1_RVT U8095 ( .A1(n8101), .A2(n8102), .Y(n8098) );
  OR2X1_RVT U8096 ( .A1(n8103), .A2(n1388), .Y(n8095) );
  AND2X1_RVT U8097 ( .A1(n8104), .A2(n8105), .Y(n8103) );
  AND2X1_RVT U8098 ( .A1(n7044), .A2(n1373), .Y(n8104) );
  OR2X1_RVT U8099 ( .A1(n83), .A2(n8106), .Y(n1373) );
  OR2X1_RVT U8100 ( .A1(n12149), .A2(n12212), .Y(n8106) );
  OR2X1_RVT U8101 ( .A1(n8107), .A2(n12191), .Y(n8094) );
  AND2X1_RVT U8102 ( .A1(n8108), .A2(n8109), .Y(n8107) );
  OR2X1_RVT U8103 ( .A1(n8110), .A2(n8055), .Y(n8109) );
  AND2X1_RVT U8104 ( .A1(n12209), .A2(n8111), .Y(n8110) );
  OR2X1_RVT U8105 ( .A1(n12189), .A2(n12185), .Y(n8111) );
  AND2X1_RVT U8106 ( .A1(n8112), .A2(n1404), .Y(n8108) );
  OR2X1_RVT U8107 ( .A1(n76), .A2(n6190), .Y(n1404) );
  OR2X1_RVT U8108 ( .A1(n8113), .A2(n1334), .Y(n8093) );
  AND4X1_RVT U8109 ( .A1(n8114), .A2(n8115), .A3(n8116), .A4(n8117), .Y(n8113)
         );
  OR2X1_RVT U8110 ( .A1(n72), .A2(n1376), .Y(n8117) );
  AND2X1_RVT U8111 ( .A1(n8118), .A2(n8119), .Y(n8116) );
  OR2X1_RVT U8112 ( .A1(n12867), .A2(n1348), .Y(n8119) );
  OR2X1_RVT U8113 ( .A1(n6198), .A2(n8120), .Y(n8118) );
  OR2X1_RVT U8114 ( .A1(n73), .A2(n12201), .Y(n8120) );
  OR2X1_RVT U8115 ( .A1(n6197), .A2(n1332), .Y(n8115) );
  OR2X1_RVT U8116 ( .A1(n12191), .A2(n8121), .Y(n8114) );
  OR2X1_RVT U8117 ( .A1(n72), .A2(n1385), .Y(n8091) );
  OR2X1_RVT U8118 ( .A1(n12204), .A2(n8122), .Y(n8090) );
  OR2X1_RVT U8119 ( .A1(n1387), .A2(n6149), .Y(n8089) );
  AND4X1_RVT U8120 ( .A1(n8123), .A2(n8124), .A3(n8125), .A4(n8126), .Y(n8045)
         );
  OR2X1_RVT U8121 ( .A1(n12871), .A2(n7033), .Y(n8126) );
  OR2X1_RVT U8122 ( .A1(n12185), .A2(n8127), .Y(n7033) );
  AND2X1_RVT U8123 ( .A1(n8128), .A2(n8129), .Y(n8125) );
  OR2X1_RVT U8124 ( .A1(n12184), .A2(n6989), .Y(n8129) );
  OR2X1_RVT U8125 ( .A1(n12870), .A2(n8130), .Y(n8128) );
  OR2X1_RVT U8126 ( .A1(n12868), .A2(n8131), .Y(n8124) );
  AND2X1_RVT U8127 ( .A1(n8132), .A2(n8133), .Y(n8123) );
  OR2X1_RVT U8128 ( .A1(n7034), .A2(n8134), .Y(n8133) );
  OR2X1_RVT U8129 ( .A1(n1312), .A2(n6159), .Y(n8132) );
  OR2X1_RVT U8130 ( .A1(n12203), .A2(n1387), .Y(n6159) );
  AND4X1_RVT U8131 ( .A1(n8136), .A2(n8137), .A3(n8138), .A4(n8139), .Y(n8135)
         );
  AND4X1_RVT U8132 ( .A1(n8140), .A2(n8141), .A3(n8142), .A4(n8143), .Y(n8139)
         );
  AND4X1_RVT U8133 ( .A1(n8144), .A2(n8145), .A3(n8146), .A4(n8147), .Y(n8143)
         );
  OR2X1_RVT U8134 ( .A1(n12339), .A2(n8149), .Y(n8142) );
  OR2X1_RVT U8135 ( .A1(n8150), .A2(n8151), .Y(n8140) );
  OR2X1_RVT U8136 ( .A1(n12768), .A2(n8152), .Y(n8151) );
  AND4X1_RVT U8137 ( .A1(n8153), .A2(n8154), .A3(n8155), .A4(n8156), .Y(n8138)
         );
  OR2X1_RVT U8138 ( .A1(n8157), .A2(n12766), .Y(n8156) );
  AND2X1_RVT U8139 ( .A1(n8158), .A2(n8159), .Y(n8157) );
  AND2X1_RVT U8140 ( .A1(n8160), .A2(n8161), .Y(n8155) );
  OR2X1_RVT U8141 ( .A1(n8162), .A2(n216), .Y(n8161) );
  AND2X1_RVT U8142 ( .A1(n8163), .A2(n8164), .Y(n8162) );
  OR2X1_RVT U8143 ( .A1(n12330), .A2(n8166), .Y(n8164) );
  OR2X1_RVT U8144 ( .A1(n8152), .A2(n8167), .Y(n8163) );
  OR2X1_RVT U8145 ( .A1(n8168), .A2(n12336), .Y(n8160) );
  AND2X1_RVT U8146 ( .A1(n8170), .A2(n8171), .Y(n8168) );
  OR2X1_RVT U8147 ( .A1(n8172), .A2(n8173), .Y(n8154) );
  AND2X1_RVT U8148 ( .A1(n8174), .A2(n8175), .Y(n8172) );
  OR2X1_RVT U8149 ( .A1(n12331), .A2(n8176), .Y(n8175) );
  AND2X1_RVT U8150 ( .A1(n8177), .A2(n8178), .Y(n8174) );
  AND2X1_RVT U8151 ( .A1(n8179), .A2(n8180), .Y(n8153) );
  OR2X1_RVT U8152 ( .A1(n8181), .A2(n12313), .Y(n8180) );
  AND2X1_RVT U8153 ( .A1(n8183), .A2(n8184), .Y(n8181) );
  OR2X1_RVT U8154 ( .A1(n8185), .A2(n8186), .Y(n8184) );
  OR2X1_RVT U8155 ( .A1(n12322), .A2(n12317), .Y(n8186) );
  OR2X1_RVT U8156 ( .A1(n8189), .A2(n8190), .Y(n8179) );
  AND2X1_RVT U8157 ( .A1(n8191), .A2(n8192), .Y(n8189) );
  AND2X1_RVT U8158 ( .A1(n8193), .A2(n8194), .Y(n8191) );
  AND4X1_RVT U8159 ( .A1(n8195), .A2(n8196), .A3(n8197), .A4(n8198), .Y(n8137)
         );
  AND4X1_RVT U8160 ( .A1(n8199), .A2(n8200), .A3(n8201), .A4(n8202), .Y(n8198)
         );
  OR2X1_RVT U8161 ( .A1(n8203), .A2(n12342), .Y(n8202) );
  AND4X1_RVT U8162 ( .A1(n8205), .A2(n8206), .A3(n8207), .A4(n8208), .Y(n8203)
         );
  OR2X1_RVT U8163 ( .A1(n8209), .A2(n8176), .Y(n8208) );
  OR2X1_RVT U8164 ( .A1(n8210), .A2(n12328), .Y(n8207) );
  OR2X1_RVT U8165 ( .A1(n8212), .A2(n12319), .Y(n8201) );
  AND4X1_RVT U8166 ( .A1(n8213), .A2(n8214), .A3(n8215), .A4(n8216), .Y(n8212)
         );
  OR2X1_RVT U8167 ( .A1(n8217), .A2(n8218), .Y(n8216) );
  OR2X1_RVT U8168 ( .A1(n12336), .A2(n12331), .Y(n8218) );
  AND2X1_RVT U8169 ( .A1(n8219), .A2(n8220), .Y(n8215) );
  OR2X1_RVT U8170 ( .A1(n12770), .A2(n8221), .Y(n8214) );
  OR2X1_RVT U8171 ( .A1(n8222), .A2(n8223), .Y(n8213) );
  AND2X1_RVT U8172 ( .A1(n8224), .A2(n8225), .Y(n8222) );
  OR2X1_RVT U8173 ( .A1(n12336), .A2(n8226), .Y(n8225) );
  OR2X1_RVT U8174 ( .A1(n8159), .A2(n8227), .Y(n8200) );
  OR2X1_RVT U8175 ( .A1(n8226), .A2(n8228), .Y(n8199) );
  OR2X1_RVT U8176 ( .A1(n8229), .A2(n8230), .Y(n8197) );
  OR2X1_RVT U8177 ( .A1(n8231), .A2(n8224), .Y(n8196) );
  OR2X1_RVT U8178 ( .A1(n8232), .A2(n8233), .Y(n8195) );
  AND4X1_RVT U8179 ( .A1(n8234), .A2(n8235), .A3(n8236), .A4(n8237), .Y(n8136)
         );
  AND2X1_RVT U8180 ( .A1(n8238), .A2(n8239), .Y(n8237) );
  OR2X1_RVT U8181 ( .A1(n8223), .A2(n8240), .Y(n8239) );
  AND2X1_RVT U8182 ( .A1(n8241), .A2(n8242), .Y(n8238) );
  OR2X1_RVT U8183 ( .A1(n8243), .A2(n8166), .Y(n8242) );
  OR2X1_RVT U8184 ( .A1(n8167), .A2(n8244), .Y(n8241) );
  OR2X1_RVT U8185 ( .A1(n214), .A2(n8245), .Y(n8236) );
  OR2X1_RVT U8186 ( .A1(n8246), .A2(n12326), .Y(n8235) );
  OR2X1_RVT U8187 ( .A1(n12329), .A2(n8248), .Y(n8234) );
  AND4X1_RVT U8188 ( .A1(n8250), .A2(n8251), .A3(n8252), .A4(n8253), .Y(n8249)
         );
  AND4X1_RVT U8189 ( .A1(n8254), .A2(n8145), .A3(n8255), .A4(n8256), .Y(n8253)
         );
  AND4X1_RVT U8190 ( .A1(n8257), .A2(n8258), .A3(n8259), .A4(n8260), .Y(n8256)
         );
  OR2X1_RVT U8191 ( .A1(n8166), .A2(n8261), .Y(n8260) );
  OR2X1_RVT U8192 ( .A1(n8262), .A2(n12341), .Y(n8261) );
  OR2X1_RVT U8193 ( .A1(n8167), .A2(n8263), .Y(n8259) );
  OR2X1_RVT U8194 ( .A1(n214), .A2(n12325), .Y(n8263) );
  OR2X1_RVT U8195 ( .A1(n8264), .A2(n8210), .Y(n8258) );
  AND2X1_RVT U8196 ( .A1(n8221), .A2(n8265), .Y(n8264) );
  OR2X1_RVT U8197 ( .A1(n8266), .A2(n8267), .Y(n8257) );
  AND2X1_RVT U8198 ( .A1(n8268), .A2(n8269), .Y(n8266) );
  AND2X1_RVT U8199 ( .A1(n8270), .A2(n8271), .Y(n8255) );
  OR2X1_RVT U8200 ( .A1(n8217), .A2(n8272), .Y(n8271) );
  OR2X1_RVT U8201 ( .A1(n8273), .A2(n12768), .Y(n8272) );
  OR2X1_RVT U8202 ( .A1(n8274), .A2(n8275), .Y(n8270) );
  OR2X1_RVT U8203 ( .A1(n8276), .A2(n12330), .Y(n8275) );
  OR2X1_RVT U8204 ( .A1(n8152), .A2(n8277), .Y(n8145) );
  AND4X1_RVT U8205 ( .A1(n8278), .A2(n8279), .A3(n8280), .A4(n8281), .Y(n8252)
         );
  AND4X1_RVT U8206 ( .A1(n8282), .A2(n8283), .A3(n8284), .A4(n8285), .Y(n8281)
         );
  OR2X1_RVT U8207 ( .A1(n8286), .A2(n12344), .Y(n8285) );
  AND2X1_RVT U8208 ( .A1(n8288), .A2(n8289), .Y(n8286) );
  OR2X1_RVT U8209 ( .A1(n12313), .A2(n8167), .Y(n8289) );
  OR2X1_RVT U8210 ( .A1(n8290), .A2(n8169), .Y(n8284) );
  AND2X1_RVT U8211 ( .A1(n8291), .A2(n8292), .Y(n8290) );
  OR2X1_RVT U8212 ( .A1(n8293), .A2(n12767), .Y(n8283) );
  AND2X1_RVT U8213 ( .A1(n8294), .A2(n8295), .Y(n8293) );
  OR2X1_RVT U8214 ( .A1(n8296), .A2(n8245), .Y(n8295) );
  AND2X1_RVT U8215 ( .A1(n12344), .A2(n12328), .Y(n8296) );
  OR2X1_RVT U8216 ( .A1(n8297), .A2(n12314), .Y(n8282) );
  AND2X1_RVT U8217 ( .A1(n8299), .A2(n8300), .Y(n8297) );
  OR2X1_RVT U8218 ( .A1(n8301), .A2(n12320), .Y(n8280) );
  AND2X1_RVT U8219 ( .A1(n8302), .A2(n8303), .Y(n8301) );
  OR2X1_RVT U8220 ( .A1(n12328), .A2(n8304), .Y(n8303) );
  AND2X1_RVT U8221 ( .A1(n8305), .A2(n8306), .Y(n8302) );
  OR2X1_RVT U8222 ( .A1(n8307), .A2(n8308), .Y(n8305) );
  OR2X1_RVT U8223 ( .A1(n8152), .A2(n8223), .Y(n8308) );
  OR2X1_RVT U8224 ( .A1(n8309), .A2(n12764), .Y(n8279) );
  AND2X1_RVT U8225 ( .A1(n8310), .A2(n8311), .Y(n8309) );
  OR2X1_RVT U8226 ( .A1(n8312), .A2(n8313), .Y(n8278) );
  AND2X1_RVT U8227 ( .A1(n8314), .A2(n8315), .Y(n8312) );
  AND2X1_RVT U8228 ( .A1(n8316), .A2(n8317), .Y(n8314) );
  OR2X1_RVT U8229 ( .A1(n216), .A2(n8245), .Y(n8317) );
  OR2X1_RVT U8230 ( .A1(n12338), .A2(n8210), .Y(n8316) );
  AND4X1_RVT U8231 ( .A1(n8318), .A2(n8319), .A3(n8320), .A4(n8321), .Y(n8251)
         );
  AND4X1_RVT U8232 ( .A1(n8322), .A2(n8323), .A3(n8324), .A4(n8325), .Y(n8321)
         );
  OR2X1_RVT U8233 ( .A1(n8245), .A2(n8244), .Y(n8325) );
  OR2X1_RVT U8234 ( .A1(n8176), .A2(n8326), .Y(n8324) );
  OR2X1_RVT U8235 ( .A1(n8209), .A2(n8327), .Y(n8323) );
  OR2X1_RVT U8236 ( .A1(n8152), .A2(n8328), .Y(n8322) );
  AND2X1_RVT U8237 ( .A1(n8329), .A2(n8330), .Y(n8320) );
  OR2X1_RVT U8238 ( .A1(n12339), .A2(n8331), .Y(n8330) );
  OR2X1_RVT U8239 ( .A1(n12318), .A2(n8228), .Y(n8329) );
  OR2X1_RVT U8240 ( .A1(n8332), .A2(n8187), .Y(n8319) );
  AND4X1_RVT U8241 ( .A1(n8333), .A2(n8334), .A3(n8335), .A4(n8336), .Y(n8332)
         );
  OR2X1_RVT U8242 ( .A1(n8337), .A2(n8152), .Y(n8335) );
  OR2X1_RVT U8243 ( .A1(n12756), .A2(n8338), .Y(n8334) );
  OR2X1_RVT U8244 ( .A1(n8339), .A2(n12764), .Y(n8333) );
  AND2X1_RVT U8245 ( .A1(n8230), .A2(n8340), .Y(n8339) );
  OR2X1_RVT U8246 ( .A1(n8232), .A2(n8341), .Y(n8318) );
  AND4X1_RVT U8247 ( .A1(n8342), .A2(n8343), .A3(n8344), .A4(n8345), .Y(n8250)
         );
  AND4X1_RVT U8248 ( .A1(n8346), .A2(n8347), .A3(n8348), .A4(n8349), .Y(n8345)
         );
  OR2X1_RVT U8249 ( .A1(n12760), .A2(n8350), .Y(n8349) );
  OR2X1_RVT U8250 ( .A1(n12761), .A2(n8351), .Y(n8348) );
  OR2X1_RVT U8251 ( .A1(n12758), .A2(n8352), .Y(n8347) );
  OR2X1_RVT U8252 ( .A1(n12312), .A2(n8353), .Y(n8346) );
  OR2X1_RVT U8253 ( .A1(n8354), .A2(n12319), .Y(n8343) );
  AND4X1_RVT U8254 ( .A1(n8356), .A2(n8357), .A3(n8358), .A4(n8359), .Y(n8355)
         );
  AND4X1_RVT U8255 ( .A1(n8360), .A2(n8361), .A3(n8362), .A4(n8363), .Y(n8359)
         );
  AND4X1_RVT U8256 ( .A1(n8364), .A2(n8141), .A3(n8311), .A4(n8365), .Y(n8363)
         );
  OR2X1_RVT U8257 ( .A1(n8366), .A2(n12755), .Y(n8141) );
  AND2X1_RVT U8258 ( .A1(n8367), .A2(n8368), .Y(n8366) );
  OR2X1_RVT U8259 ( .A1(n8185), .A2(n8369), .Y(n8368) );
  OR2X1_RVT U8260 ( .A1(n8370), .A2(n8267), .Y(n8367) );
  OR2X1_RVT U8261 ( .A1(n8371), .A2(n8226), .Y(n8364) );
  AND2X1_RVT U8262 ( .A1(n8372), .A2(n8373), .Y(n8371) );
  OR2X1_RVT U8263 ( .A1(n12760), .A2(n8210), .Y(n8373) );
  OR2X1_RVT U8264 ( .A1(n8374), .A2(n8169), .Y(n8362) );
  AND2X1_RVT U8265 ( .A1(n8375), .A2(n8376), .Y(n8374) );
  OR2X1_RVT U8266 ( .A1(n8377), .A2(n12766), .Y(n8376) );
  AND2X1_RVT U8267 ( .A1(n8217), .A2(n8378), .Y(n8377) );
  OR2X1_RVT U8268 ( .A1(n8379), .A2(n12339), .Y(n8361) );
  AND2X1_RVT U8269 ( .A1(n8380), .A2(n8381), .Y(n8379) );
  OR2X1_RVT U8270 ( .A1(n8210), .A2(n8176), .Y(n8381) );
  OR2X1_RVT U8271 ( .A1(n8382), .A2(n12322), .Y(n8360) );
  AND2X1_RVT U8272 ( .A1(n8294), .A2(n8383), .Y(n8382) );
  OR2X1_RVT U8273 ( .A1(n8223), .A2(n8384), .Y(n8294) );
  AND4X1_RVT U8274 ( .A1(n8385), .A2(n8386), .A3(n8387), .A4(n8388), .Y(n8358)
         );
  OR2X1_RVT U8275 ( .A1(n8389), .A2(n12329), .Y(n8388) );
  AND2X1_RVT U8276 ( .A1(n8390), .A2(n8391), .Y(n8389) );
  OR2X1_RVT U8277 ( .A1(n8267), .A2(n8167), .Y(n8391) );
  AND2X1_RVT U8278 ( .A1(n8392), .A2(n8393), .Y(n8390) );
  OR2X1_RVT U8279 ( .A1(n8307), .A2(n8369), .Y(n8392) );
  AND2X1_RVT U8280 ( .A1(n8394), .A2(n8395), .Y(n8387) );
  OR2X1_RVT U8281 ( .A1(n8396), .A2(n8298), .Y(n8395) );
  AND2X1_RVT U8282 ( .A1(n8397), .A2(n8206), .Y(n8396) );
  OR2X1_RVT U8283 ( .A1(n8152), .A2(n8267), .Y(n8206) );
  OR2X1_RVT U8284 ( .A1(n8398), .A2(n216), .Y(n8394) );
  AND2X1_RVT U8285 ( .A1(n8399), .A2(n8400), .Y(n8398) );
  OR2X1_RVT U8286 ( .A1(n8401), .A2(n12331), .Y(n8400) );
  AND2X1_RVT U8287 ( .A1(n8402), .A2(n8403), .Y(n8401) );
  OR2X1_RVT U8288 ( .A1(n12326), .A2(n8217), .Y(n8403) );
  OR2X1_RVT U8289 ( .A1(n12770), .A2(n12328), .Y(n8402) );
  AND2X1_RVT U8290 ( .A1(n8268), .A2(n8378), .Y(n8399) );
  OR2X1_RVT U8291 ( .A1(n8298), .A2(n8404), .Y(n8268) );
  OR2X1_RVT U8292 ( .A1(n12765), .A2(n12761), .Y(n8404) );
  OR2X1_RVT U8293 ( .A1(n8405), .A2(n8287), .Y(n8386) );
  AND4X1_RVT U8294 ( .A1(n8246), .A2(n8406), .A3(n8407), .A4(n8408), .Y(n8405)
         );
  OR2X1_RVT U8295 ( .A1(n12330), .A2(n8267), .Y(n8408) );
  AND2X1_RVT U8296 ( .A1(n8409), .A2(n8410), .Y(n8407) );
  OR2X1_RVT U8297 ( .A1(n12770), .A2(n12339), .Y(n8406) );
  AND2X1_RVT U8298 ( .A1(n8411), .A2(n8412), .Y(n8246) );
  OR2X1_RVT U8299 ( .A1(n8413), .A2(n214), .Y(n8412) );
  OR2X1_RVT U8300 ( .A1(n8210), .A2(n12755), .Y(n8411) );
  AND2X1_RVT U8301 ( .A1(n8414), .A2(n8415), .Y(n8385) );
  OR2X1_RVT U8302 ( .A1(n8416), .A2(n12757), .Y(n8415) );
  AND2X1_RVT U8303 ( .A1(n8417), .A2(n8418), .Y(n8416) );
  OR2X1_RVT U8304 ( .A1(n8419), .A2(n12333), .Y(n8418) );
  AND2X1_RVT U8305 ( .A1(n8420), .A2(n8421), .Y(n8419) );
  AND2X1_RVT U8306 ( .A1(n8422), .A2(n8423), .Y(n8417) );
  OR2X1_RVT U8307 ( .A1(n8424), .A2(n12342), .Y(n8414) );
  AND4X1_RVT U8308 ( .A1(n8425), .A2(n8426), .A3(n8427), .A4(n8428), .Y(n8424)
         );
  OR2X1_RVT U8309 ( .A1(n12769), .A2(n8429), .Y(n8427) );
  OR2X1_RVT U8310 ( .A1(n214), .A2(n8224), .Y(n8426) );
  OR2X1_RVT U8311 ( .A1(n8313), .A2(n8267), .Y(n8425) );
  AND4X1_RVT U8312 ( .A1(n8430), .A2(n8431), .A3(n8432), .A4(n8433), .Y(n8357)
         );
  AND2X1_RVT U8313 ( .A1(n8434), .A2(n8277), .Y(n8433) );
  OR2X1_RVT U8314 ( .A1(n12317), .A2(n8243), .Y(n8277) );
  AND2X1_RVT U8315 ( .A1(n8435), .A2(n8436), .Y(n8434) );
  OR2X1_RVT U8316 ( .A1(n8437), .A2(n8192), .Y(n8436) );
  OR2X1_RVT U8317 ( .A1(n8244), .A2(n8304), .Y(n8435) );
  OR2X1_RVT U8318 ( .A1(n214), .A2(n8438), .Y(n8432) );
  OR2X1_RVT U8319 ( .A1(n12768), .A2(n8439), .Y(n8431) );
  OR2X1_RVT U8320 ( .A1(n8313), .A2(n8440), .Y(n8430) );
  AND4X1_RVT U8321 ( .A1(n8441), .A2(n8442), .A3(n8443), .A4(n8444), .Y(n8356)
         );
  AND2X1_RVT U8322 ( .A1(n8445), .A2(n8446), .Y(n8444) );
  OR2X1_RVT U8323 ( .A1(n12312), .A2(n8447), .Y(n8446) );
  AND2X1_RVT U8324 ( .A1(n8448), .A2(n8449), .Y(n8445) );
  OR2X1_RVT U8325 ( .A1(n8209), .A2(n8219), .Y(n8449) );
  OR2X1_RVT U8326 ( .A1(n12333), .A2(n8269), .Y(n8219) );
  OR2X1_RVT U8327 ( .A1(n12319), .A2(n8450), .Y(n8448) );
  OR2X1_RVT U8328 ( .A1(n8190), .A2(n8183), .Y(n8443) );
  OR2X1_RVT U8329 ( .A1(n8276), .A2(n8451), .Y(n8183) );
  OR2X1_RVT U8330 ( .A1(n12764), .A2(n8452), .Y(n8442) );
  OR2X1_RVT U8331 ( .A1(n12331), .A2(n8310), .Y(n8441) );
  OR2X1_RVT U8332 ( .A1(n12755), .A2(n8372), .Y(n8310) );
  AND4X1_RVT U8333 ( .A1(n8454), .A2(n8455), .A3(n8456), .A4(n8457), .Y(n8453)
         );
  AND4X1_RVT U8334 ( .A1(n8458), .A2(n8459), .A3(n8460), .A4(n8461), .Y(n8457)
         );
  OR2X1_RVT U8335 ( .A1(n224), .A2(n8462), .Y(n8461) );
  OR2X1_RVT U8336 ( .A1(n8463), .A2(n12344), .Y(n8462) );
  AND2X1_RVT U8337 ( .A1(n12333), .A2(n8229), .Y(n8463) );
  AND2X1_RVT U8338 ( .A1(n8144), .A2(n8464), .Y(n8460) );
  OR2X1_RVT U8339 ( .A1(n12322), .A2(n8465), .Y(n8144) );
  OR2X1_RVT U8340 ( .A1(n224), .A2(n8223), .Y(n8465) );
  OR2X1_RVT U8341 ( .A1(n8466), .A2(n8152), .Y(n8459) );
  AND2X1_RVT U8342 ( .A1(n8467), .A2(n8468), .Y(n8466) );
  AND2X1_RVT U8343 ( .A1(n8469), .A2(n8470), .Y(n8458) );
  OR2X1_RVT U8344 ( .A1(n8471), .A2(n8472), .Y(n8470) );
  AND2X1_RVT U8345 ( .A1(n8473), .A2(n8233), .Y(n8471) );
  OR2X1_RVT U8346 ( .A1(n8474), .A2(n8224), .Y(n8469) );
  AND2X1_RVT U8347 ( .A1(n8409), .A2(n8243), .Y(n8474) );
  OR2X1_RVT U8348 ( .A1(n12320), .A2(n8475), .Y(n8409) );
  OR2X1_RVT U8349 ( .A1(n12770), .A2(n12330), .Y(n8475) );
  AND4X1_RVT U8350 ( .A1(n8476), .A2(n8477), .A3(n8478), .A4(n8479), .Y(n8456)
         );
  OR2X1_RVT U8351 ( .A1(n8480), .A2(n12760), .Y(n8479) );
  AND2X1_RVT U8352 ( .A1(n8292), .A2(n8481), .Y(n8480) );
  OR2X1_RVT U8353 ( .A1(n12768), .A2(n8337), .Y(n8292) );
  AND2X1_RVT U8354 ( .A1(n8482), .A2(n8483), .Y(n8478) );
  OR2X1_RVT U8355 ( .A1(n8484), .A2(n12758), .Y(n8483) );
  AND2X1_RVT U8356 ( .A1(n8485), .A2(n8486), .Y(n8484) );
  OR2X1_RVT U8357 ( .A1(n8187), .A2(n8429), .Y(n8486) );
  OR2X1_RVT U8358 ( .A1(n8487), .A2(n12756), .Y(n8482) );
  AND2X1_RVT U8359 ( .A1(n8488), .A2(n8489), .Y(n8487) );
  OR2X1_RVT U8360 ( .A1(n8490), .A2(n12333), .Y(n8477) );
  AND2X1_RVT U8361 ( .A1(n8491), .A2(n8492), .Y(n8490) );
  AND2X1_RVT U8362 ( .A1(n8493), .A2(n8494), .Y(n8491) );
  AND2X1_RVT U8363 ( .A1(n8495), .A2(n8496), .Y(n8476) );
  OR2X1_RVT U8364 ( .A1(n8497), .A2(n8413), .Y(n8496) );
  AND2X1_RVT U8365 ( .A1(n8498), .A2(n8244), .Y(n8497) );
  AND2X1_RVT U8366 ( .A1(n8499), .A2(n8500), .Y(n8498) );
  OR2X1_RVT U8367 ( .A1(n8501), .A2(n12336), .Y(n8495) );
  AND2X1_RVT U8368 ( .A1(n8502), .A2(n8503), .Y(n8501) );
  OR2X1_RVT U8369 ( .A1(n12767), .A2(n12338), .Y(n8503) );
  AND2X1_RVT U8370 ( .A1(n8233), .A2(n8504), .Y(n8502) );
  AND4X1_RVT U8371 ( .A1(n8505), .A2(n8506), .A3(n8507), .A4(n8508), .Y(n8455)
         );
  AND2X1_RVT U8372 ( .A1(n8509), .A2(n8510), .Y(n8508) );
  OR2X1_RVT U8373 ( .A1(n8226), .A2(n8300), .Y(n8510) );
  OR2X1_RVT U8374 ( .A1(n12762), .A2(n8233), .Y(n8300) );
  AND2X1_RVT U8375 ( .A1(n8511), .A2(n8512), .Y(n8509) );
  OR2X1_RVT U8376 ( .A1(n8378), .A2(n8192), .Y(n8512) );
  OR2X1_RVT U8377 ( .A1(n12769), .A2(n12329), .Y(n8192) );
  OR2X1_RVT U8378 ( .A1(n8276), .A2(n8326), .Y(n8511) );
  OR2X1_RVT U8379 ( .A1(n12757), .A2(n8513), .Y(n8326) );
  OR2X1_RVT U8380 ( .A1(n8514), .A2(n12312), .Y(n8507) );
  AND4X1_RVT U8381 ( .A1(n8515), .A2(n8516), .A3(n8517), .A4(n8518), .Y(n8514)
         );
  OR2X1_RVT U8382 ( .A1(n8451), .A2(n8224), .Y(n8517) );
  OR2X1_RVT U8383 ( .A1(n8519), .A2(n8221), .Y(n8516) );
  OR2X1_RVT U8384 ( .A1(n12766), .A2(n8176), .Y(n8515) );
  OR2X1_RVT U8385 ( .A1(n8520), .A2(n12313), .Y(n8506) );
  AND2X1_RVT U8386 ( .A1(n8521), .A2(n8522), .Y(n8520) );
  OR2X1_RVT U8387 ( .A1(n8451), .A2(n8176), .Y(n8522) );
  AND2X1_RVT U8388 ( .A1(n8523), .A2(n8452), .Y(n8521) );
  OR2X1_RVT U8389 ( .A1(n8224), .A2(n8524), .Y(n8452) );
  OR2X1_RVT U8390 ( .A1(n12757), .A2(n12769), .Y(n8524) );
  OR2X1_RVT U8391 ( .A1(n8525), .A2(n12320), .Y(n8505) );
  AND4X1_RVT U8392 ( .A1(n8526), .A2(n8439), .A3(n8248), .A4(n8220), .Y(n8525)
         );
  OR2X1_RVT U8393 ( .A1(n8245), .A2(n8527), .Y(n8220) );
  OR2X1_RVT U8394 ( .A1(n12759), .A2(n8182), .Y(n8527) );
  OR2X1_RVT U8395 ( .A1(n8307), .A2(n8341), .Y(n8248) );
  OR2X1_RVT U8396 ( .A1(n8226), .A2(n8528), .Y(n8439) );
  OR2X1_RVT U8397 ( .A1(n12344), .A2(n12313), .Y(n8528) );
  OR2X1_RVT U8398 ( .A1(n8185), .A2(n8529), .Y(n8526) );
  OR2X1_RVT U8399 ( .A1(n8530), .A2(n12318), .Y(n8529) );
  AND4X1_RVT U8400 ( .A1(n8531), .A2(n8532), .A3(n8533), .A4(n8534), .Y(n8454)
         );
  AND2X1_RVT U8401 ( .A1(n8535), .A2(n8536), .Y(n8534) );
  AND2X1_RVT U8402 ( .A1(n8537), .A2(n8538), .Y(n8535) );
  OR2X1_RVT U8403 ( .A1(n8217), .A2(n8492), .Y(n8538) );
  OR2X1_RVT U8404 ( .A1(n8229), .A2(n8539), .Y(n8492) );
  OR2X1_RVT U8405 ( .A1(n12758), .A2(n12760), .Y(n8539) );
  OR2X1_RVT U8406 ( .A1(n12765), .A2(n8540), .Y(n8537) );
  OR2X1_RVT U8407 ( .A1(n12329), .A2(n8541), .Y(n8533) );
  OR2X1_RVT U8408 ( .A1(n12768), .A2(n8542), .Y(n8532) );
  OR2X1_RVT U8409 ( .A1(n8229), .A2(n8543), .Y(n8531) );
  AND4X1_RVT U8410 ( .A1(n8545), .A2(n8546), .A3(n8547), .A4(n8548), .Y(n8544)
         );
  AND4X1_RVT U8411 ( .A1(n8549), .A2(n8550), .A3(n8551), .A4(n8552), .Y(n8548)
         );
  AND4X1_RVT U8412 ( .A1(n8553), .A2(n8554), .A3(n8146), .A4(n8555), .Y(n8552)
         );
  OR2X1_RVT U8413 ( .A1(n8287), .A2(n8556), .Y(n8146) );
  OR2X1_RVT U8414 ( .A1(n8378), .A2(n216), .Y(n8556) );
  OR2X1_RVT U8415 ( .A1(n8150), .A2(n8557), .Y(n8554) );
  OR2X1_RVT U8416 ( .A1(n12763), .A2(n12766), .Y(n8557) );
  OR2X1_RVT U8417 ( .A1(n8413), .A2(n8558), .Y(n8553) );
  OR2X1_RVT U8418 ( .A1(n8559), .A2(n8187), .Y(n8558) );
  AND2X1_RVT U8419 ( .A1(n12333), .A2(n8287), .Y(n8559) );
  OR2X1_RVT U8420 ( .A1(n8560), .A2(n12339), .Y(n8551) );
  AND2X1_RVT U8421 ( .A1(n8428), .A2(n8500), .Y(n8560) );
  OR2X1_RVT U8422 ( .A1(n216), .A2(n8561), .Y(n8500) );
  OR2X1_RVT U8423 ( .A1(n12312), .A2(n12762), .Y(n8561) );
  OR2X1_RVT U8424 ( .A1(n8217), .A2(n8562), .Y(n8428) );
  OR2X1_RVT U8425 ( .A1(n12760), .A2(n8209), .Y(n8562) );
  OR2X1_RVT U8426 ( .A1(n8563), .A2(n8167), .Y(n8550) );
  AND2X1_RVT U8427 ( .A1(n8564), .A2(n8372), .Y(n8563) );
  OR2X1_RVT U8428 ( .A1(n8273), .A2(n8267), .Y(n8549) );
  AND4X1_RVT U8429 ( .A1(n8565), .A2(n8566), .A3(n8567), .A4(n8568), .Y(n8547)
         );
  AND2X1_RVT U8430 ( .A1(n8569), .A2(n8570), .Y(n8568) );
  OR2X1_RVT U8431 ( .A1(n8571), .A2(n12333), .Y(n8570) );
  AND2X1_RVT U8432 ( .A1(n8572), .A2(n8240), .Y(n8571) );
  AND2X1_RVT U8433 ( .A1(n8573), .A2(n8574), .Y(n8569) );
  OR2X1_RVT U8434 ( .A1(n8575), .A2(n8223), .Y(n8574) );
  AND2X1_RVT U8435 ( .A1(n8194), .A2(n8166), .Y(n8575) );
  OR2X1_RVT U8436 ( .A1(n12768), .A2(n8265), .Y(n8194) );
  OR2X1_RVT U8437 ( .A1(n8576), .A2(n8276), .Y(n8573) );
  AND2X1_RVT U8438 ( .A1(n8468), .A2(n8577), .Y(n8576) );
  OR2X1_RVT U8439 ( .A1(n12769), .A2(n8304), .Y(n8468) );
  OR2X1_RVT U8440 ( .A1(n8578), .A2(n12760), .Y(n8567) );
  AND2X1_RVT U8441 ( .A1(n8171), .A2(n8579), .Y(n8578) );
  OR2X1_RVT U8442 ( .A1(n8307), .A2(n8231), .Y(n8579) );
  OR2X1_RVT U8443 ( .A1(n8210), .A2(n8413), .Y(n8171) );
  OR2X1_RVT U8444 ( .A1(n8580), .A2(n214), .Y(n8566) );
  AND2X1_RVT U8445 ( .A1(n8221), .A2(n8581), .Y(n8580) );
  OR2X1_RVT U8446 ( .A1(n8582), .A2(n12317), .Y(n8581) );
  AND2X1_RVT U8447 ( .A1(n8583), .A2(n8584), .Y(n8582) );
  OR2X1_RVT U8448 ( .A1(n12761), .A2(n8204), .Y(n8584) );
  OR2X1_RVT U8449 ( .A1(n12344), .A2(n8307), .Y(n8221) );
  OR2X1_RVT U8450 ( .A1(n8585), .A2(n8291), .Y(n8565) );
  AND2X1_RVT U8451 ( .A1(n8224), .A2(n8269), .Y(n8585) );
  OR2X1_RVT U8452 ( .A1(n12757), .A2(n8152), .Y(n8269) );
  AND4X1_RVT U8453 ( .A1(n8586), .A2(n8587), .A3(n8588), .A4(n8589), .Y(n8546)
         );
  AND4X1_RVT U8454 ( .A1(n8590), .A2(n8591), .A3(n8592), .A4(n8593), .Y(n8589)
         );
  OR2X1_RVT U8455 ( .A1(n8594), .A2(n12768), .Y(n8593) );
  AND2X1_RVT U8456 ( .A1(n8327), .A2(n8595), .Y(n8594) );
  OR2X1_RVT U8457 ( .A1(n12341), .A2(n8176), .Y(n8595) );
  OR2X1_RVT U8458 ( .A1(n8596), .A2(n8169), .Y(n8592) );
  AND2X1_RVT U8459 ( .A1(n8597), .A2(n8598), .Y(n8596) );
  OR2X1_RVT U8460 ( .A1(n8599), .A2(n8204), .Y(n8598) );
  AND2X1_RVT U8461 ( .A1(n8229), .A2(n8217), .Y(n8599) );
  AND2X1_RVT U8462 ( .A1(n8231), .A2(n8473), .Y(n8597) );
  OR2X1_RVT U8463 ( .A1(n12342), .A2(n8369), .Y(n8473) );
  OR2X1_RVT U8464 ( .A1(n8600), .A2(n12331), .Y(n8591) );
  AND2X1_RVT U8465 ( .A1(n8601), .A2(n8602), .Y(n8600) );
  OR2X1_RVT U8466 ( .A1(n8217), .A2(n8603), .Y(n8602) );
  AND2X1_RVT U8467 ( .A1(n8299), .A2(n8493), .Y(n8601) );
  OR2X1_RVT U8468 ( .A1(n8209), .A2(n8384), .Y(n8493) );
  OR2X1_RVT U8469 ( .A1(n8182), .A2(n8604), .Y(n8299) );
  OR2X1_RVT U8470 ( .A1(n8605), .A2(n8152), .Y(n8590) );
  AND4X1_RVT U8471 ( .A1(n8606), .A2(n8607), .A3(n8608), .A4(n8541), .Y(n8605)
         );
  OR2X1_RVT U8472 ( .A1(n8245), .A2(n8609), .Y(n8541) );
  OR2X1_RVT U8473 ( .A1(n12312), .A2(n8209), .Y(n8609) );
  OR2X1_RVT U8474 ( .A1(n12765), .A2(n8451), .Y(n8607) );
  OR2X1_RVT U8475 ( .A1(n8210), .A2(n8307), .Y(n8606) );
  OR2X1_RVT U8476 ( .A1(n8378), .A2(n8420), .Y(n8588) );
  OR2X1_RVT U8477 ( .A1(n8610), .A2(n12315), .Y(n8587) );
  AND4X1_RVT U8478 ( .A1(n8611), .A2(n8612), .A3(n8254), .A4(n8352), .Y(n8610)
         );
  OR2X1_RVT U8479 ( .A1(n8176), .A2(n8341), .Y(n8352) );
  OR2X1_RVT U8480 ( .A1(n12765), .A2(n214), .Y(n8341) );
  OR2X1_RVT U8481 ( .A1(n8169), .A2(n8233), .Y(n8254) );
  OR2X1_RVT U8482 ( .A1(n12757), .A2(n8604), .Y(n8586) );
  AND4X1_RVT U8483 ( .A1(n8613), .A2(n8614), .A3(n8615), .A4(n8616), .Y(n8545)
         );
  OR2X1_RVT U8484 ( .A1(n12320), .A2(n8617), .Y(n8616) );
  AND2X1_RVT U8485 ( .A1(n8618), .A2(n8619), .Y(n8615) );
  OR2X1_RVT U8486 ( .A1(n12341), .A2(n8372), .Y(n8619) );
  OR2X1_RVT U8487 ( .A1(n8159), .A2(n8233), .Y(n8618) );
  OR2X1_RVT U8488 ( .A1(n216), .A2(n8190), .Y(n8233) );
  OR2X1_RVT U8489 ( .A1(n12344), .A2(n8351), .Y(n8614) );
  OR2X1_RVT U8490 ( .A1(n8226), .A2(n8620), .Y(n8351) );
  AND2X1_RVT U8491 ( .A1(n8621), .A2(n8622), .Y(n8613) );
  OR2X1_RVT U8492 ( .A1(n12313), .A2(n8623), .Y(n8622) );
  OR2X1_RVT U8493 ( .A1(n8229), .A2(n8178), .Y(n8621) );
  OR2X1_RVT U8494 ( .A1(n8152), .A2(n8437), .Y(n8178) );
  AND4X1_RVT U8495 ( .A1(n8625), .A2(n8626), .A3(n8627), .A4(n8628), .Y(n8624)
         );
  AND4X1_RVT U8496 ( .A1(n8629), .A2(n8630), .A3(n8631), .A4(n8632), .Y(n8628)
         );
  AND4X1_RVT U8497 ( .A1(n8365), .A2(n8555), .A3(n8633), .A4(n8634), .Y(n8632)
         );
  OR2X1_RVT U8498 ( .A1(n8635), .A2(n8636), .Y(n8555) );
  OR2X1_RVT U8499 ( .A1(n8150), .A2(n8420), .Y(n8365) );
  OR2X1_RVT U8500 ( .A1(n12766), .A2(n12329), .Y(n8420) );
  AND4X1_RVT U8501 ( .A1(n8623), .A2(n8489), .A3(n8612), .A4(n8147), .Y(n8631)
         );
  OR2X1_RVT U8502 ( .A1(n8637), .A2(n8337), .Y(n8147) );
  OR2X1_RVT U8503 ( .A1(n8152), .A2(n8638), .Y(n8612) );
  OR2X1_RVT U8504 ( .A1(n8185), .A2(n214), .Y(n8489) );
  OR2X1_RVT U8505 ( .A1(n8176), .A2(n8639), .Y(n8623) );
  OR2X1_RVT U8506 ( .A1(n12319), .A2(n12339), .Y(n8639) );
  AND4X1_RVT U8507 ( .A1(n8640), .A2(n8641), .A3(n8642), .A4(n8643), .Y(n8630)
         );
  OR2X1_RVT U8508 ( .A1(n8429), .A2(n8644), .Y(n8643) );
  OR2X1_RVT U8509 ( .A1(n12339), .A2(n8209), .Y(n8644) );
  OR2X1_RVT U8510 ( .A1(n8338), .A2(n8645), .Y(n8642) );
  OR2X1_RVT U8511 ( .A1(n12767), .A2(n8226), .Y(n8645) );
  OR2X1_RVT U8512 ( .A1(n8564), .A2(n8646), .Y(n8641) );
  OR2X1_RVT U8513 ( .A1(n8647), .A2(n8223), .Y(n8646) );
  OR2X1_RVT U8514 ( .A1(n12336), .A2(n8648), .Y(n8640) );
  OR2X1_RVT U8515 ( .A1(n8649), .A2(n12319), .Y(n8648) );
  AND2X1_RVT U8516 ( .A1(n8437), .A2(n8650), .Y(n8649) );
  AND2X1_RVT U8517 ( .A1(n8651), .A2(n8652), .Y(n8629) );
  OR2X1_RVT U8518 ( .A1(n8653), .A2(n8204), .Y(n8652) );
  AND2X1_RVT U8519 ( .A1(n8654), .A2(n8655), .Y(n8653) );
  OR2X1_RVT U8520 ( .A1(n12318), .A2(n8397), .Y(n8655) );
  OR2X1_RVT U8521 ( .A1(n12322), .A2(n8472), .Y(n8654) );
  AND2X1_RVT U8522 ( .A1(n8656), .A2(n8657), .Y(n8651) );
  OR2X1_RVT U8523 ( .A1(n8658), .A2(n8243), .Y(n8657) );
  AND2X1_RVT U8524 ( .A1(n8659), .A2(n8660), .Y(n8658) );
  OR2X1_RVT U8525 ( .A1(n12325), .A2(n224), .Y(n8660) );
  NAND2X1_RVT U8526 ( .A1(n8226), .A2(n12759), .Y(n8659) );
  OR2X1_RVT U8527 ( .A1(n8661), .A2(n216), .Y(n8656) );
  AND2X1_RVT U8528 ( .A1(n8450), .A2(n8327), .Y(n8661) );
  OR2X1_RVT U8529 ( .A1(n8176), .A2(n8662), .Y(n8327) );
  OR2X1_RVT U8530 ( .A1(n12770), .A2(n12314), .Y(n8662) );
  AND4X1_RVT U8531 ( .A1(n8344), .A2(n8663), .A3(n8536), .A4(n8664), .Y(n8627)
         );
  AND4X1_RVT U8532 ( .A1(n8665), .A2(n8666), .A3(n8667), .A4(n8668), .Y(n8664)
         );
  OR2X1_RVT U8533 ( .A1(n8307), .A2(n8228), .Y(n8668) );
  OR2X1_RVT U8534 ( .A1(n8245), .A2(n8274), .Y(n8667) );
  OR2X1_RVT U8535 ( .A1(n12758), .A2(n8499), .Y(n8666) );
  OR2X1_RVT U8536 ( .A1(n8223), .A2(n8205), .Y(n8499) );
  OR2X1_RVT U8537 ( .A1(n12766), .A2(n8287), .Y(n8205) );
  OR2X1_RVT U8538 ( .A1(n12328), .A2(n8328), .Y(n8665) );
  OR2X1_RVT U8539 ( .A1(n8209), .A2(n8437), .Y(n8328) );
  OR2X1_RVT U8540 ( .A1(n12312), .A2(n8413), .Y(n8437) );
  AND2X1_RVT U8541 ( .A1(n8669), .A2(n8670), .Y(n8536) );
  OR2X1_RVT U8542 ( .A1(n8671), .A2(n8276), .Y(n8670) );
  OR2X1_RVT U8543 ( .A1(n12338), .A2(n216), .Y(n8671) );
  OR2X1_RVT U8544 ( .A1(n8672), .A2(n8159), .Y(n8669) );
  OR2X1_RVT U8545 ( .A1(n12757), .A2(n8276), .Y(n8159) );
  OR2X1_RVT U8546 ( .A1(n8173), .A2(n8223), .Y(n8672) );
  OR2X1_RVT U8547 ( .A1(n12320), .A2(n8542), .Y(n8663) );
  AND2X1_RVT U8548 ( .A1(n8673), .A2(n8674), .Y(n8344) );
  OR2X1_RVT U8549 ( .A1(n8227), .A2(n8265), .Y(n8674) );
  OR2X1_RVT U8550 ( .A1(n8675), .A2(n8676), .Y(n8673) );
  AND4X1_RVT U8551 ( .A1(n8677), .A2(n8678), .A3(n8679), .A4(n8680), .Y(n8626)
         );
  OR2X1_RVT U8552 ( .A1(n8681), .A2(n8413), .Y(n8680) );
  AND2X1_RVT U8553 ( .A1(n8682), .A2(n8422), .Y(n8681) );
  OR2X1_RVT U8554 ( .A1(n12326), .A2(n8638), .Y(n8422) );
  OR2X1_RVT U8555 ( .A1(n8683), .A2(n12763), .Y(n8679) );
  AND2X1_RVT U8556 ( .A1(n8350), .A2(n8315), .Y(n8683) );
  OR2X1_RVT U8557 ( .A1(n12757), .A2(n8291), .Y(n8315) );
  OR2X1_RVT U8558 ( .A1(n8684), .A2(n8370), .Y(n8678) );
  AND2X1_RVT U8559 ( .A1(n8685), .A2(n8686), .Y(n8684) );
  OR2X1_RVT U8560 ( .A1(n12315), .A2(n8229), .Y(n8686) );
  AND2X1_RVT U8561 ( .A1(n8687), .A2(n8267), .Y(n8685) );
  OR2X1_RVT U8562 ( .A1(n214), .A2(n8226), .Y(n8687) );
  OR2X1_RVT U8563 ( .A1(n8688), .A2(n8167), .Y(n8677) );
  AND2X1_RVT U8564 ( .A1(n8689), .A2(n8690), .Y(n8688) );
  NAND2X1_RVT U8565 ( .A1(n8152), .A2(n8530), .Y(n8690) );
  AND2X1_RVT U8566 ( .A1(n8691), .A2(n8380), .Y(n8689) );
  OR2X1_RVT U8567 ( .A1(n8313), .A2(n8638), .Y(n8380) );
  OR2X1_RVT U8568 ( .A1(n12335), .A2(n8692), .Y(n8691) );
  AND4X1_RVT U8569 ( .A1(n8693), .A2(n8694), .A3(n8695), .A4(n8696), .Y(n8625)
         );
  OR2X1_RVT U8570 ( .A1(n8697), .A2(n8190), .Y(n8696) );
  AND2X1_RVT U8571 ( .A1(n8698), .A2(n8331), .Y(n8697) );
  AND2X1_RVT U8572 ( .A1(n8699), .A2(n8353), .Y(n8698) );
  OR2X1_RVT U8573 ( .A1(n216), .A2(n8676), .Y(n8353) );
  OR2X1_RVT U8574 ( .A1(n12314), .A2(n8287), .Y(n8676) );
  OR2X1_RVT U8575 ( .A1(n8700), .A2(n12331), .Y(n8695) );
  AND2X1_RVT U8576 ( .A1(n8701), .A2(n8702), .Y(n8700) );
  OR2X1_RVT U8577 ( .A1(n8703), .A2(n12755), .Y(n8702) );
  AND2X1_RVT U8578 ( .A1(n8704), .A2(n8705), .Y(n8703) );
  OR2X1_RVT U8579 ( .A1(n12313), .A2(n8564), .Y(n8705) );
  OR2X1_RVT U8580 ( .A1(n12762), .A2(n8210), .Y(n8704) );
  AND2X1_RVT U8581 ( .A1(n8706), .A2(n8707), .Y(n8701) );
  OR2X1_RVT U8582 ( .A1(n8176), .A2(n8708), .Y(n8706) );
  OR2X1_RVT U8583 ( .A1(n8709), .A2(n8210), .Y(n8694) );
  AND4X1_RVT U8584 ( .A1(n8710), .A2(n8711), .A3(n8712), .A4(n8176), .Y(n8709)
         );
  OR2X1_RVT U8585 ( .A1(n12763), .A2(n8226), .Y(n8712) );
  OR2X1_RVT U8586 ( .A1(n12325), .A2(n8245), .Y(n8711) );
  OR2X1_RVT U8587 ( .A1(n8298), .A2(n8276), .Y(n8710) );
  OR2X1_RVT U8588 ( .A1(n8713), .A2(n8152), .Y(n8693) );
  AND4X1_RVT U8589 ( .A1(n8577), .A2(n8714), .A3(n8375), .A4(n8291), .Y(n8713)
         );
  OR2X1_RVT U8590 ( .A1(n8245), .A2(n8708), .Y(n8375) );
  OR2X1_RVT U8591 ( .A1(n8413), .A2(n8620), .Y(n8714) );
  OR2X1_RVT U8592 ( .A1(n12319), .A2(n8378), .Y(n8577) );
  AND4X1_RVT U8593 ( .A1(n8716), .A2(n8717), .A3(n8718), .A4(n8719), .Y(n8715)
         );
  AND4X1_RVT U8594 ( .A1(n8228), .A2(n8464), .A3(n8720), .A4(n8721), .Y(n8719)
         );
  AND4X1_RVT U8595 ( .A1(n8543), .A2(n8488), .A3(n8633), .A4(n8634), .Y(n8721)
         );
  OR2X1_RVT U8596 ( .A1(n8636), .A2(n8149), .Y(n8634) );
  OR2X1_RVT U8597 ( .A1(n12761), .A2(n8267), .Y(n8149) );
  OR2X1_RVT U8598 ( .A1(n8166), .A2(n8675), .Y(n8633) );
  OR2X1_RVT U8599 ( .A1(n12766), .A2(n12333), .Y(n8675) );
  OR2X1_RVT U8600 ( .A1(n12755), .A2(n8287), .Y(n8166) );
  OR2X1_RVT U8601 ( .A1(n12767), .A2(n8185), .Y(n8488) );
  OR2X1_RVT U8602 ( .A1(n12342), .A2(n12326), .Y(n8185) );
  OR2X1_RVT U8603 ( .A1(n8307), .A2(n8722), .Y(n8543) );
  OR2X1_RVT U8604 ( .A1(n12333), .A2(n8211), .Y(n8722) );
  OR2X1_RVT U8605 ( .A1(n8209), .A2(n8723), .Y(n8720) );
  OR2X1_RVT U8606 ( .A1(n8337), .A2(n12324), .Y(n8723) );
  OR2X1_RVT U8607 ( .A1(n8276), .A2(n8724), .Y(n8464) );
  OR2X1_RVT U8608 ( .A1(n8210), .A2(n12331), .Y(n8724) );
  OR2X1_RVT U8609 ( .A1(n12759), .A2(n8635), .Y(n8228) );
  OR2X1_RVT U8610 ( .A1(n12326), .A2(n8227), .Y(n8635) );
  AND4X1_RVT U8611 ( .A1(n8725), .A2(n8726), .A3(n8727), .A4(n8728), .Y(n8718)
         );
  AND4X1_RVT U8612 ( .A1(n8729), .A2(n8730), .A3(n8731), .A4(n8732), .Y(n8728)
         );
  OR2X1_RVT U8613 ( .A1(n8243), .A2(n8733), .Y(n8732) );
  OR2X1_RVT U8614 ( .A1(n12315), .A2(n8313), .Y(n8733) );
  OR2X1_RVT U8615 ( .A1(n8226), .A2(n8734), .Y(n8731) );
  OR2X1_RVT U8616 ( .A1(n8735), .A2(n8190), .Y(n8734) );
  AND2X1_RVT U8617 ( .A1(n8169), .A2(n8229), .Y(n8735) );
  OR2X1_RVT U8618 ( .A1(n8736), .A2(n8737), .Y(n8730) );
  AND2X1_RVT U8619 ( .A1(n8384), .A2(n8340), .Y(n8736) );
  OR2X1_RVT U8620 ( .A1(n12760), .A2(n224), .Y(n8340) );
  OR2X1_RVT U8621 ( .A1(n12756), .A2(n12336), .Y(n8384) );
  OR2X1_RVT U8622 ( .A1(n8738), .A2(n8224), .Y(n8729) );
  AND2X1_RVT U8623 ( .A1(n8620), .A2(n8739), .Y(n8738) );
  OR2X1_RVT U8624 ( .A1(n12758), .A2(n216), .Y(n8739) );
  OR2X1_RVT U8625 ( .A1(n8740), .A2(n12338), .Y(n8727) );
  AND2X1_RVT U8626 ( .A1(n8611), .A2(n8741), .Y(n8740) );
  OR2X1_RVT U8627 ( .A1(n8217), .A2(n8564), .Y(n8741) );
  OR2X1_RVT U8628 ( .A1(n12319), .A2(n8429), .Y(n8611) );
  OR2X1_RVT U8629 ( .A1(n12762), .A2(n8217), .Y(n8429) );
  OR2X1_RVT U8630 ( .A1(n8742), .A2(n8378), .Y(n8726) );
  AND2X1_RVT U8631 ( .A1(n8331), .A2(n8603), .Y(n8742) );
  OR2X1_RVT U8632 ( .A1(n8187), .A2(n8276), .Y(n8331) );
  OR2X1_RVT U8633 ( .A1(n8743), .A2(n8267), .Y(n8725) );
  AND2X1_RVT U8634 ( .A1(n8230), .A2(n8232), .Y(n8743) );
  AND4X1_RVT U8635 ( .A1(n8744), .A2(n8745), .A3(n8746), .A4(n8747), .Y(n8717)
         );
  AND4X1_RVT U8636 ( .A1(n8748), .A2(n8749), .A3(n8750), .A4(n8751), .Y(n8747)
         );
  OR2X1_RVT U8637 ( .A1(n8752), .A2(n12322), .Y(n8751) );
  AND2X1_RVT U8638 ( .A1(n8158), .A2(n8450), .Y(n8752) );
  OR2X1_RVT U8639 ( .A1(n8307), .A2(n8338), .Y(n8450) );
  OR2X1_RVT U8640 ( .A1(n12325), .A2(n8190), .Y(n8338) );
  OR2X1_RVT U8641 ( .A1(n12329), .A2(n8753), .Y(n8158) );
  OR2X1_RVT U8642 ( .A1(n12312), .A2(n12318), .Y(n8753) );
  OR2X1_RVT U8643 ( .A1(n8754), .A2(n12336), .Y(n8750) );
  AND2X1_RVT U8644 ( .A1(n8467), .A2(n8755), .Y(n8754) );
  OR2X1_RVT U8645 ( .A1(n12341), .A2(n214), .Y(n8755) );
  OR2X1_RVT U8646 ( .A1(n12339), .A2(n8274), .Y(n8467) );
  OR2X1_RVT U8647 ( .A1(n8756), .A2(n12317), .Y(n8749) );
  AND2X1_RVT U8648 ( .A1(n8485), .A2(n8757), .Y(n8756) );
  OR2X1_RVT U8649 ( .A1(n12342), .A2(n8210), .Y(n8757) );
  OR2X1_RVT U8650 ( .A1(n8152), .A2(n8758), .Y(n8485) );
  OR2X1_RVT U8651 ( .A1(n8759), .A2(n8211), .Y(n8748) );
  AND2X1_RVT U8652 ( .A1(n8760), .A2(n8761), .Y(n8759) );
  OR2X1_RVT U8653 ( .A1(n8267), .A2(n12339), .Y(n8761) );
  AND2X1_RVT U8654 ( .A1(n8762), .A2(n8243), .Y(n8760) );
  OR2X1_RVT U8655 ( .A1(n8229), .A2(n8190), .Y(n8243) );
  OR2X1_RVT U8656 ( .A1(n12314), .A2(n8274), .Y(n8762) );
  OR2X1_RVT U8657 ( .A1(n12770), .A2(n8229), .Y(n8274) );
  OR2X1_RVT U8658 ( .A1(n8763), .A2(n8287), .Y(n8746) );
  AND4X1_RVT U8659 ( .A1(n8764), .A2(n8765), .A3(n8440), .A4(n8350), .Y(n8763)
         );
  OR2X1_RVT U8660 ( .A1(n8413), .A2(n8513), .Y(n8350) );
  OR2X1_RVT U8661 ( .A1(n8245), .A2(n8692), .Y(n8440) );
  OR2X1_RVT U8662 ( .A1(n12320), .A2(n12313), .Y(n8692) );
  OR2X1_RVT U8663 ( .A1(n216), .A2(n8167), .Y(n8765) );
  OR2X1_RVT U8664 ( .A1(n214), .A2(n12339), .Y(n8764) );
  OR2X1_RVT U8665 ( .A1(n8766), .A2(n8223), .Y(n8745) );
  AND2X1_RVT U8666 ( .A1(n8767), .A2(n8244), .Y(n8766) );
  AND2X1_RVT U8667 ( .A1(n8699), .A2(n8494), .Y(n8767) );
  OR2X1_RVT U8668 ( .A1(n8768), .A2(n12767), .Y(n8494) );
  AND2X1_RVT U8669 ( .A1(n8265), .A2(n8769), .Y(n8768) );
  OR2X1_RVT U8670 ( .A1(n12317), .A2(n8152), .Y(n8769) );
  OR2X1_RVT U8671 ( .A1(n8313), .A2(n8451), .Y(n8699) );
  OR2X1_RVT U8672 ( .A1(n8298), .A2(n8187), .Y(n8451) );
  OR2X1_RVT U8673 ( .A1(n8770), .A2(n8291), .Y(n8744) );
  AND2X1_RVT U8674 ( .A1(n8771), .A2(n12325), .Y(n8770) );
  AND2X1_RVT U8675 ( .A1(n8772), .A2(n8472), .Y(n8771) );
  OR2X1_RVT U8676 ( .A1(n8313), .A2(n8413), .Y(n8772) );
  AND4X1_RVT U8677 ( .A1(n8773), .A2(n8774), .A3(n8775), .A4(n8776), .Y(n8716)
         );
  AND2X1_RVT U8678 ( .A1(n8777), .A2(n8778), .Y(n8776) );
  OR2X1_RVT U8679 ( .A1(n12763), .A2(n8393), .Y(n8778) );
  OR2X1_RVT U8680 ( .A1(n12333), .A2(n8779), .Y(n8393) );
  OR2X1_RVT U8681 ( .A1(n8209), .A2(n8298), .Y(n8779) );
  AND2X1_RVT U8682 ( .A1(n8780), .A2(n8781), .Y(n8777) );
  OR2X1_RVT U8683 ( .A1(n8182), .A2(n8193), .Y(n8781) );
  OR2X1_RVT U8684 ( .A1(n8226), .A2(n8421), .Y(n8193) );
  OR2X1_RVT U8685 ( .A1(n12759), .A2(n8187), .Y(n8421) );
  OR2X1_RVT U8686 ( .A1(n8229), .A2(n8306), .Y(n8780) );
  OR2X1_RVT U8687 ( .A1(n8217), .A2(n8782), .Y(n8306) );
  OR2X1_RVT U8688 ( .A1(n8217), .A2(n8397), .Y(n8775) );
  OR2X1_RVT U8689 ( .A1(n216), .A2(n12335), .Y(n8397) );
  OR2X1_RVT U8690 ( .A1(n8783), .A2(n8173), .Y(n8774) );
  AND4X1_RVT U8691 ( .A1(n8784), .A2(n8785), .A3(n8786), .A4(n8787), .Y(n8783)
         );
  OR2X1_RVT U8692 ( .A1(n12757), .A2(n8788), .Y(n8786) );
  OR2X1_RVT U8693 ( .A1(n8789), .A2(n12764), .Y(n8788) );
  AND2X1_RVT U8694 ( .A1(n8224), .A2(n8790), .Y(n8789) );
  OR2X1_RVT U8695 ( .A1(n12328), .A2(n8791), .Y(n8785) );
  OR2X1_RVT U8696 ( .A1(n8530), .A2(n8167), .Y(n8791) );
  OR2X1_RVT U8697 ( .A1(n8150), .A2(n8176), .Y(n8784) );
  OR2X1_RVT U8698 ( .A1(n12761), .A2(n8276), .Y(n8176) );
  OR2X1_RVT U8699 ( .A1(n8650), .A2(n8564), .Y(n8773) );
  OR2X1_RVT U8700 ( .A1(n12344), .A2(n8187), .Y(n8564) );
  AND4X1_RVT U8701 ( .A1(n8793), .A2(n8794), .A3(n8795), .A4(n8796), .Y(n8792)
         );
  AND4X1_RVT U8702 ( .A1(n8797), .A2(n8798), .A3(n8799), .A4(n8800), .Y(n8796)
         );
  AND4X1_RVT U8703 ( .A1(n8801), .A2(n8802), .A3(n8803), .A4(n8804), .Y(n8800)
         );
  OR2X1_RVT U8704 ( .A1(n8638), .A2(n8782), .Y(n8804) );
  OR2X1_RVT U8705 ( .A1(n12760), .A2(n12338), .Y(n8782) );
  OR2X1_RVT U8706 ( .A1(n12312), .A2(n12322), .Y(n8638) );
  OR2X1_RVT U8707 ( .A1(n8805), .A2(n8224), .Y(n8803) );
  AND2X1_RVT U8708 ( .A1(n8170), .A2(n8737), .Y(n8805) );
  OR2X1_RVT U8709 ( .A1(n216), .A2(n8806), .Y(n8170) );
  OR2X1_RVT U8710 ( .A1(n12312), .A2(n12757), .Y(n8806) );
  OR2X1_RVT U8711 ( .A1(n8807), .A2(n8152), .Y(n8802) );
  OR2X1_RVT U8712 ( .A1(n12326), .A2(n8313), .Y(n8152) );
  AND2X1_RVT U8713 ( .A1(n8288), .A2(n8808), .Y(n8807) );
  OR2X1_RVT U8714 ( .A1(n8167), .A2(n8369), .Y(n8808) );
  OR2X1_RVT U8715 ( .A1(n12330), .A2(n12318), .Y(n8167) );
  OR2X1_RVT U8716 ( .A1(n8413), .A2(n8809), .Y(n8288) );
  OR2X1_RVT U8717 ( .A1(n12768), .A2(n12333), .Y(n8809) );
  OR2X1_RVT U8718 ( .A1(n8810), .A2(n8211), .Y(n8801) );
  AND2X1_RVT U8719 ( .A1(n8608), .A2(n8811), .Y(n8810) );
  OR2X1_RVT U8720 ( .A1(n8812), .A2(n12757), .Y(n8811) );
  AND2X1_RVT U8721 ( .A1(n8267), .A2(n8620), .Y(n8812) );
  OR2X1_RVT U8722 ( .A1(n12765), .A2(n8229), .Y(n8620) );
  OR2X1_RVT U8723 ( .A1(n12339), .A2(n8813), .Y(n8608) );
  OR2X1_RVT U8724 ( .A1(n12770), .A2(n12766), .Y(n8813) );
  OR2X1_RVT U8725 ( .A1(n8814), .A2(n12317), .Y(n8799) );
  AND2X1_RVT U8726 ( .A1(n8815), .A2(n8816), .Y(n8814) );
  OR2X1_RVT U8727 ( .A1(n8817), .A2(n8313), .Y(n8816) );
  AND2X1_RVT U8728 ( .A1(n8378), .A2(n8818), .Y(n8817) );
  OR2X1_RVT U8729 ( .A1(n8169), .A2(n8291), .Y(n8815) );
  OR2X1_RVT U8730 ( .A1(n12331), .A2(n8227), .Y(n8291) );
  OR2X1_RVT U8731 ( .A1(n8819), .A2(n12766), .Y(n8798) );
  AND2X1_RVT U8732 ( .A1(n8383), .A2(n8542), .Y(n8819) );
  OR2X1_RVT U8733 ( .A1(n12329), .A2(n8820), .Y(n8542) );
  OR2X1_RVT U8734 ( .A1(n8223), .A2(n12318), .Y(n8820) );
  OR2X1_RVT U8735 ( .A1(n8169), .A2(n8650), .Y(n8383) );
  OR2X1_RVT U8736 ( .A1(n12318), .A2(n12333), .Y(n8650) );
  OR2X1_RVT U8737 ( .A1(n8821), .A2(n12315), .Y(n8797) );
  AND2X1_RVT U8738 ( .A1(n8423), .A2(n8822), .Y(n8821) );
  OR2X1_RVT U8739 ( .A1(n8637), .A2(n8217), .Y(n8822) );
  OR2X1_RVT U8740 ( .A1(n8276), .A2(n8758), .Y(n8423) );
  OR2X1_RVT U8741 ( .A1(n12765), .A2(n216), .Y(n8758) );
  AND2X1_RVT U8742 ( .A1(n12319), .A2(n12768), .Y(n8519) );
  AND4X1_RVT U8743 ( .A1(n8823), .A2(n8824), .A3(n8825), .A4(n8826), .Y(n8795)
         );
  AND4X1_RVT U8744 ( .A1(n8827), .A2(n8828), .A3(n8829), .A4(n8830), .Y(n8826)
         );
  OR2X1_RVT U8745 ( .A1(n8831), .A2(n12324), .Y(n8830) );
  AND2X1_RVT U8746 ( .A1(n8410), .A2(n8481), .Y(n8831) );
  OR2X1_RVT U8747 ( .A1(n8226), .A2(n8737), .Y(n8481) );
  OR2X1_RVT U8748 ( .A1(n12768), .A2(n8223), .Y(n8737) );
  OR2X1_RVT U8749 ( .A1(n12755), .A2(n12314), .Y(n8226) );
  OR2X1_RVT U8750 ( .A1(n12315), .A2(n8513), .Y(n8410) );
  OR2X1_RVT U8751 ( .A1(n12319), .A2(n12333), .Y(n8513) );
  OR2X1_RVT U8752 ( .A1(n8832), .A2(n12764), .Y(n8829) );
  AND2X1_RVT U8753 ( .A1(n8572), .A2(n8833), .Y(n8832) );
  OR2X1_RVT U8754 ( .A1(n8530), .A2(n8240), .Y(n8833) );
  OR2X1_RVT U8755 ( .A1(n8413), .A2(n8834), .Y(n8240) );
  OR2X1_RVT U8756 ( .A1(n12344), .A2(n12320), .Y(n8834) );
  OR2X1_RVT U8757 ( .A1(n12328), .A2(n8835), .Y(n8572) );
  OR2X1_RVT U8758 ( .A1(n8413), .A2(n8209), .Y(n8835) );
  OR2X1_RVT U8759 ( .A1(n8836), .A2(n12770), .Y(n8828) );
  AND2X1_RVT U8760 ( .A1(n8518), .A2(n8447), .Y(n8836) );
  OR2X1_RVT U8761 ( .A1(n8229), .A2(n8265), .Y(n8447) );
  OR2X1_RVT U8762 ( .A1(n12762), .A2(n8413), .Y(n8265) );
  OR2X1_RVT U8763 ( .A1(n8637), .A2(n8245), .Y(n8518) );
  OR2X1_RVT U8764 ( .A1(n12325), .A2(n12767), .Y(n8637) );
  OR2X1_RVT U8765 ( .A1(n8837), .A2(n8287), .Y(n8827) );
  AND2X1_RVT U8766 ( .A1(n8838), .A2(n8839), .Y(n8837) );
  OR2X1_RVT U8767 ( .A1(n8209), .A2(n8636), .Y(n8839) );
  OR2X1_RVT U8768 ( .A1(n12764), .A2(n224), .Y(n8636) );
  AND2X1_RVT U8769 ( .A1(n8840), .A2(n8504), .Y(n8838) );
  OR2X1_RVT U8770 ( .A1(n8217), .A2(n8841), .Y(n8504) );
  OR2X1_RVT U8771 ( .A1(n12341), .A2(n12320), .Y(n8841) );
  OR2X1_RVT U8772 ( .A1(n8273), .A2(n8210), .Y(n8825) );
  OR2X1_RVT U8773 ( .A1(n12757), .A2(n8169), .Y(n8273) );
  OR2X1_RVT U8774 ( .A1(n8842), .A2(n8173), .Y(n8824) );
  AND2X1_RVT U8775 ( .A1(n8843), .A2(n8354), .Y(n8842) );
  AND2X1_RVT U8776 ( .A1(n8844), .A2(n8845), .Y(n8354) );
  OR2X1_RVT U8777 ( .A1(n12329), .A2(n8378), .Y(n8845) );
  OR2X1_RVT U8778 ( .A1(n8276), .A2(n8150), .Y(n8844) );
  OR2X1_RVT U8779 ( .A1(n12314), .A2(n8223), .Y(n8150) );
  AND2X1_RVT U8780 ( .A1(n8846), .A2(n8540), .Y(n8843) );
  OR2X1_RVT U8781 ( .A1(n8307), .A2(n8790), .Y(n8540) );
  OR2X1_RVT U8782 ( .A1(n12759), .A2(n214), .Y(n8790) );
  OR2X1_RVT U8783 ( .A1(n8169), .A2(n8336), .Y(n8846) );
  OR2X1_RVT U8784 ( .A1(n12313), .A2(n8847), .Y(n8336) );
  OR2X1_RVT U8785 ( .A1(n12755), .A2(n12342), .Y(n8847) );
  OR2X1_RVT U8786 ( .A1(n8848), .A2(n12755), .Y(n8823) );
  AND4X1_RVT U8787 ( .A1(n8849), .A2(n8850), .A3(n8851), .A4(n8682), .Y(n8848)
         );
  OR2X1_RVT U8788 ( .A1(n8223), .A2(n8603), .Y(n8682) );
  OR2X1_RVT U8789 ( .A1(n12760), .A2(n12766), .Y(n8603) );
  OR2X1_RVT U8790 ( .A1(n8223), .A2(n8852), .Y(n8851) );
  OR2X1_RVT U8791 ( .A1(n12319), .A2(n12324), .Y(n8852) );
  OR2X1_RVT U8792 ( .A1(n12765), .A2(n8182), .Y(n8223) );
  OR2X1_RVT U8793 ( .A1(n8853), .A2(n8304), .Y(n8850) );
  OR2X1_RVT U8794 ( .A1(n12313), .A2(n8148), .Y(n8304) );
  AND2X1_RVT U8795 ( .A1(n8287), .A2(n8854), .Y(n8853) );
  OR2X1_RVT U8796 ( .A1(n12763), .A2(n8187), .Y(n8854) );
  OR2X1_RVT U8797 ( .A1(n12759), .A2(n12324), .Y(n8287) );
  OR2X1_RVT U8798 ( .A1(n12761), .A2(n8818), .Y(n8849) );
  OR2X1_RVT U8799 ( .A1(n12765), .A2(n8227), .Y(n8818) );
  OR2X1_RVT U8800 ( .A1(n8173), .A2(n214), .Y(n8227) );
  AND4X1_RVT U8801 ( .A1(n8855), .A2(n8856), .A3(n8857), .A4(n8858), .Y(n8794)
         );
  AND4X1_RVT U8802 ( .A1(n8859), .A2(n8860), .A3(n8861), .A4(n8862), .Y(n8858)
         );
  OR2X1_RVT U8803 ( .A1(n8245), .A2(n8372), .Y(n8862) );
  OR2X1_RVT U8804 ( .A1(n12326), .A2(n8267), .Y(n8372) );
  OR2X1_RVT U8805 ( .A1(n12330), .A2(n8413), .Y(n8245) );
  OR2X1_RVT U8806 ( .A1(n8232), .A2(n8708), .Y(n8861) );
  OR2X1_RVT U8807 ( .A1(n12769), .A2(n12313), .Y(n8708) );
  OR2X1_RVT U8808 ( .A1(n8298), .A2(n8224), .Y(n8232) );
  OR2X1_RVT U8809 ( .A1(n8217), .A2(n8244), .Y(n8860) );
  OR2X1_RVT U8810 ( .A1(n12322), .A2(n12335), .Y(n8244) );
  OR2X1_RVT U8811 ( .A1(n12312), .A2(n12756), .Y(n8217) );
  OR2X1_RVT U8812 ( .A1(n224), .A2(n8583), .Y(n8859) );
  OR2X1_RVT U8813 ( .A1(n12320), .A2(n8370), .Y(n8583) );
  OR2X1_RVT U8814 ( .A1(n8187), .A2(n8617), .Y(n8857) );
  OR2X1_RVT U8815 ( .A1(n224), .A2(n8863), .Y(n8617) );
  OR2X1_RVT U8816 ( .A1(n12762), .A2(n12333), .Y(n8863) );
  AND2X1_RVT U8817 ( .A1(n12314), .A2(n12317), .Y(n8647) );
  OR2X1_RVT U8818 ( .A1(n8229), .A2(n8177), .Y(n8856) );
  OR2X1_RVT U8819 ( .A1(n12342), .A2(n8864), .Y(n8177) );
  OR2X1_RVT U8820 ( .A1(n12763), .A2(n12755), .Y(n8864) );
  OR2X1_RVT U8821 ( .A1(n12319), .A2(n8209), .Y(n8229) );
  OR2X1_RVT U8822 ( .A1(n8276), .A2(n8840), .Y(n8855) );
  OR2X1_RVT U8823 ( .A1(n12315), .A2(n8231), .Y(n8840) );
  OR2X1_RVT U8824 ( .A1(n12765), .A2(n12766), .Y(n8231) );
  AND4X1_RVT U8825 ( .A1(n8865), .A2(n8342), .A3(n8866), .A4(n8867), .Y(n8793)
         );
  OR2X1_RVT U8826 ( .A1(n12319), .A2(n8787), .Y(n8867) );
  OR2X1_RVT U8827 ( .A1(n12761), .A2(n8337), .Y(n8787) );
  OR2X1_RVT U8828 ( .A1(n12317), .A2(n8378), .Y(n8337) );
  OR2X1_RVT U8829 ( .A1(n12312), .A2(n8204), .Y(n8378) );
  AND2X1_RVT U8830 ( .A1(n8868), .A2(n8869), .Y(n8866) );
  OR2X1_RVT U8831 ( .A1(n12341), .A2(n8707), .Y(n8869) );
  OR2X1_RVT U8832 ( .A1(n8276), .A2(n8369), .Y(n8707) );
  OR2X1_RVT U8833 ( .A1(n12319), .A2(n12313), .Y(n8369) );
  OR2X1_RVT U8834 ( .A1(n12314), .A2(n8165), .Y(n8204) );
  OR2X1_RVT U8835 ( .A1(n12768), .A2(n8438), .Y(n8868) );
  OR2X1_RVT U8836 ( .A1(n12338), .A2(n8472), .Y(n8438) );
  OR2X1_RVT U8837 ( .A1(n12760), .A2(n12755), .Y(n8472) );
  OR2X1_RVT U8838 ( .A1(n12758), .A2(n12330), .Y(n8148) );
  AND2X1_RVT U8839 ( .A1(n8870), .A2(n8871), .Y(n8342) );
  OR2X1_RVT U8840 ( .A1(n8224), .A2(n8210), .Y(n8871) );
  OR2X1_RVT U8841 ( .A1(n12767), .A2(n8182), .Y(n8210) );
  AND2X1_RVT U8842 ( .A1(n8209), .A2(n8173), .Y(n8262) );
  OR2X1_RVT U8843 ( .A1(n12325), .A2(n8276), .Y(n8224) );
  OR2X1_RVT U8844 ( .A1(n12756), .A2(n8313), .Y(n8276) );
  OR2X1_RVT U8845 ( .A1(n8872), .A2(n8267), .Y(n8870) );
  OR2X1_RVT U8846 ( .A1(n12319), .A2(n214), .Y(n8267) );
  AND2X1_RVT U8847 ( .A1(n12769), .A2(n12312), .Y(n8530) );
  OR2X1_RVT U8848 ( .A1(n12318), .A2(n8370), .Y(n8872) );
  OR2X1_RVT U8849 ( .A1(n12765), .A2(n12335), .Y(n8370) );
  AND2X1_RVT U8850 ( .A1(n8873), .A2(n8874), .Y(n8865) );
  OR2X1_RVT U8851 ( .A1(n8190), .A2(n8523), .Y(n8874) );
  OR2X1_RVT U8852 ( .A1(n12320), .A2(n8230), .Y(n8523) );
  OR2X1_RVT U8853 ( .A1(n12335), .A2(n8307), .Y(n8230) );
  OR2X1_RVT U8854 ( .A1(n12315), .A2(n12318), .Y(n8307) );
  OR2X1_RVT U8855 ( .A1(n12762), .A2(n12760), .Y(n8169) );
  OR2X1_RVT U8856 ( .A1(n12770), .A2(n12764), .Y(n8190) );
  XOR2X1_RVT U8857 ( .A1(key[44]), .A2(state[44]), .Y(n8165) );
  OR2X1_RVT U8858 ( .A1(n8182), .A2(n8311), .Y(n8873) );
  OR2X1_RVT U8859 ( .A1(n8413), .A2(n8604), .Y(n8311) );
  OR2X1_RVT U8860 ( .A1(n12322), .A2(n8211), .Y(n8604) );
  OR2X1_RVT U8861 ( .A1(n12763), .A2(n8313), .Y(n8211) );
  XOR2X1_RVT U8862 ( .A1(key[42]), .A2(state[42]), .Y(n8313) );
  XOR2X1_RVT U8863 ( .A1(key[43]), .A2(state[43]), .Y(n8247) );
  OR2X1_RVT U8864 ( .A1(n12768), .A2(n12320), .Y(n8187) );
  XOR2X1_RVT U8865 ( .A1(key[45]), .A2(state[45]), .Y(n8173) );
  XOR2X1_RVT U8866 ( .A1(key[46]), .A2(state[46]), .Y(n8209) );
  OR2X1_RVT U8867 ( .A1(n12758), .A2(n12318), .Y(n8413) );
  XOR2X1_RVT U8868 ( .A1(key[40]), .A2(state[40]), .Y(n8188) );
  XOR2X1_RVT U8869 ( .A1(key[41]), .A2(state[41]), .Y(n8298) );
  XOR2X1_RVT U8870 ( .A1(key[47]), .A2(state[47]), .Y(n8182) );
  AND4X1_RVT U8871 ( .A1(n8876), .A2(n8877), .A3(n8878), .A4(n8879), .Y(n8875)
         );
  AND4X1_RVT U8872 ( .A1(n8880), .A2(n8881), .A3(n8882), .A4(n8883), .Y(n8879)
         );
  AND4X1_RVT U8873 ( .A1(n8884), .A2(n8885), .A3(n8886), .A4(n8887), .Y(n8883)
         );
  OR2X1_RVT U8874 ( .A1(n6176), .A2(n8888), .Y(n8886) );
  OR2X1_RVT U8875 ( .A1(n8889), .A2(n12189), .Y(n8888) );
  AND2X1_RVT U8876 ( .A1(n69), .A2(n12876), .Y(n8889) );
  OR2X1_RVT U8877 ( .A1(n1342), .A2(n8890), .Y(n8885) );
  OR2X1_RVT U8878 ( .A1(n8891), .A2(n12926), .Y(n8884) );
  AND2X1_RVT U8879 ( .A1(n8892), .A2(n8893), .Y(n8891) );
  OR2X1_RVT U8880 ( .A1(n8894), .A2(n69), .Y(n8893) );
  AND2X1_RVT U8881 ( .A1(n83), .A2(n8895), .Y(n8894) );
  OR2X1_RVT U8882 ( .A1(n8063), .A2(n1350), .Y(n8895) );
  OR2X1_RVT U8883 ( .A1(n8896), .A2(n73), .Y(n8882) );
  AND2X1_RVT U8884 ( .A1(n1372), .A2(n8897), .Y(n8896) );
  OR2X1_RVT U8885 ( .A1(n1325), .A2(n7007), .Y(n8897) );
  OR2X1_RVT U8886 ( .A1(n1332), .A2(n8898), .Y(n1372) );
  OR2X1_RVT U8887 ( .A1(n12149), .A2(n12201), .Y(n8898) );
  OR2X1_RVT U8888 ( .A1(n8899), .A2(n12204), .Y(n8881) );
  AND2X1_RVT U8889 ( .A1(n1313), .A2(n8900), .Y(n8899) );
  OR2X1_RVT U8890 ( .A1(n8901), .A2(n6143), .Y(n8900) );
  OR2X1_RVT U8891 ( .A1(n12199), .A2(n78), .Y(n1313) );
  OR2X1_RVT U8892 ( .A1(n8902), .A2(n12875), .Y(n8880) );
  AND2X1_RVT U8893 ( .A1(n1374), .A2(n8903), .Y(n8902) );
  OR2X1_RVT U8894 ( .A1(n8904), .A2(n12149), .Y(n8903) );
  AND2X1_RVT U8895 ( .A1(n6973), .A2(n8905), .Y(n8904) );
  OR2X1_RVT U8896 ( .A1(n1325), .A2(n6198), .Y(n8905) );
  OR2X1_RVT U8897 ( .A1(n12203), .A2(n1332), .Y(n6973) );
  OR2X1_RVT U8898 ( .A1(n12204), .A2(n1347), .Y(n1374) );
  AND4X1_RVT U8899 ( .A1(n8906), .A2(n8907), .A3(n8908), .A4(n8909), .Y(n8878)
         );
  OR2X1_RVT U8900 ( .A1(n8910), .A2(n1356), .Y(n8909) );
  AND2X1_RVT U8901 ( .A1(n8911), .A2(n8912), .Y(n8910) );
  AND2X1_RVT U8902 ( .A1(n6975), .A2(n1301), .Y(n8911) );
  OR2X1_RVT U8903 ( .A1(n12194), .A2(n7013), .Y(n1301) );
  OR2X1_RVT U8904 ( .A1(n12150), .A2(n8127), .Y(n6975) );
  AND2X1_RVT U8905 ( .A1(n8913), .A2(n8914), .Y(n8908) );
  OR2X1_RVT U8906 ( .A1(n8915), .A2(n71), .Y(n8914) );
  AND2X1_RVT U8907 ( .A1(n6976), .A2(n8916), .Y(n8915) );
  OR2X1_RVT U8908 ( .A1(n72), .A2(n8917), .Y(n8916) );
  OR2X1_RVT U8909 ( .A1(n78), .A2(n6180), .Y(n6976) );
  OR2X1_RVT U8910 ( .A1(n8918), .A2(n8919), .Y(n8913) );
  AND2X1_RVT U8911 ( .A1(n8920), .A2(n8921), .Y(n8918) );
  OR2X1_RVT U8912 ( .A1(n12198), .A2(n8922), .Y(n8921) );
  NAND2X1_RVT U8913 ( .A1(n1307), .A2(n12185), .Y(n8922) );
  AND2X1_RVT U8914 ( .A1(n8923), .A2(n8105), .Y(n8920) );
  OR2X1_RVT U8915 ( .A1(n78), .A2(n8924), .Y(n8105) );
  OR2X1_RVT U8916 ( .A1(n8917), .A2(n8925), .Y(n8907) );
  AND2X1_RVT U8917 ( .A1(n8926), .A2(n8927), .Y(n8906) );
  OR2X1_RVT U8918 ( .A1(n8928), .A2(n12194), .Y(n8927) );
  AND2X1_RVT U8919 ( .A1(n8929), .A2(n8930), .Y(n8928) );
  OR2X1_RVT U8920 ( .A1(n6128), .A2(n8931), .Y(n8930) );
  OR2X1_RVT U8921 ( .A1(n1361), .A2(n12188), .Y(n8931) );
  AND2X1_RVT U8922 ( .A1(n8083), .A2(n6158), .Y(n8929) );
  OR2X1_RVT U8923 ( .A1(n6198), .A2(n8932), .Y(n6158) );
  OR2X1_RVT U8924 ( .A1(n12199), .A2(n8933), .Y(n8083) );
  OR2X1_RVT U8925 ( .A1(n1325), .A2(n12186), .Y(n8933) );
  OR2X1_RVT U8926 ( .A1(n8934), .A2(n12869), .Y(n8926) );
  AND4X1_RVT U8927 ( .A1(n6149), .A2(n8935), .A3(n70), .A4(n8936), .Y(n8934)
         );
  AND4X1_RVT U8928 ( .A1(n8937), .A2(n8131), .A3(n7045), .A4(n6191), .Y(n8936)
         );
  OR2X1_RVT U8929 ( .A1(n8919), .A2(n7030), .Y(n6191) );
  OR2X1_RVT U8930 ( .A1(n12184), .A2(n6184), .Y(n7045) );
  OR2X1_RVT U8931 ( .A1(n1300), .A2(n6172), .Y(n8131) );
  OR2X1_RVT U8932 ( .A1(n12211), .A2(n12875), .Y(n6149) );
  AND4X1_RVT U8933 ( .A1(n8938), .A2(n8939), .A3(n8940), .A4(n8941), .Y(n8877)
         );
  AND2X1_RVT U8934 ( .A1(n8942), .A2(n8943), .Y(n8941) );
  OR2X1_RVT U8935 ( .A1(n1387), .A2(n6192), .Y(n8943) );
  OR2X1_RVT U8936 ( .A1(n12192), .A2(n78), .Y(n1387) );
  AND2X1_RVT U8937 ( .A1(n8944), .A2(n8945), .Y(n8942) );
  OR2X1_RVT U8938 ( .A1(n6143), .A2(n7008), .Y(n8945) );
  OR2X1_RVT U8939 ( .A1(n6139), .A2(n8946), .Y(n8944) );
  OR2X1_RVT U8940 ( .A1(n1325), .A2(n8947), .Y(n8940) );
  OR2X1_RVT U8941 ( .A1(n6132), .A2(n8121), .Y(n8939) );
  OR2X1_RVT U8942 ( .A1(n85), .A2(n6967), .Y(n8938) );
  OR2X1_RVT U8943 ( .A1(n1314), .A2(n8121), .Y(n6967) );
  AND4X1_RVT U8944 ( .A1(n8948), .A2(n8949), .A3(n8950), .A4(n6206), .Y(n8876)
         );
  OR2X1_RVT U8945 ( .A1(n78), .A2(n8951), .Y(n6206) );
  OR2X1_RVT U8946 ( .A1(n12206), .A2(n6972), .Y(n8951) );
  OR2X1_RVT U8947 ( .A1(n85), .A2(n7034), .Y(n6972) );
  AND2X1_RVT U8948 ( .A1(n8952), .A2(n8953), .Y(n8950) );
  OR2X1_RVT U8949 ( .A1(n76), .A2(n8954), .Y(n8953) );
  OR2X1_RVT U8950 ( .A1(n8063), .A2(n7019), .Y(n8952) );
  OR2X1_RVT U8951 ( .A1(n12209), .A2(n6184), .Y(n7019) );
  OR2X1_RVT U8952 ( .A1(n73), .A2(n12211), .Y(n6184) );
  OR2X1_RVT U8953 ( .A1(n12872), .A2(n8955), .Y(n8949) );
  AND2X1_RVT U8954 ( .A1(n8956), .A2(n8957), .Y(n8948) );
  OR2X1_RVT U8955 ( .A1(n1391), .A2(n7005), .Y(n8957) );
  OR2X1_RVT U8956 ( .A1(n1341), .A2(n1397), .Y(n8956) );
  OR2X1_RVT U8957 ( .A1(n6145), .A2(n8958), .Y(n1397) );
  OR2X1_RVT U8958 ( .A1(n12874), .A2(n7034), .Y(n8958) );
  AND4X1_RVT U8959 ( .A1(n8960), .A2(n8961), .A3(n8962), .A4(n8963), .Y(n8959)
         );
  AND4X1_RVT U8960 ( .A1(n8964), .A2(n8965), .A3(n8966), .A4(n8967), .Y(n8963)
         );
  AND4X1_RVT U8961 ( .A1(n8968), .A2(n8969), .A3(n8970), .A4(n8971), .Y(n8967)
         );
  OR2X1_RVT U8962 ( .A1(n12306), .A2(n8973), .Y(n8966) );
  OR2X1_RVT U8963 ( .A1(n8974), .A2(n8975), .Y(n8964) );
  OR2X1_RVT U8964 ( .A1(n12752), .A2(n8976), .Y(n8975) );
  AND4X1_RVT U8965 ( .A1(n8977), .A2(n8978), .A3(n8979), .A4(n8980), .Y(n8962)
         );
  OR2X1_RVT U8966 ( .A1(n8981), .A2(n12750), .Y(n8980) );
  AND2X1_RVT U8967 ( .A1(n8982), .A2(n8983), .Y(n8981) );
  AND2X1_RVT U8968 ( .A1(n8984), .A2(n8985), .Y(n8979) );
  OR2X1_RVT U8969 ( .A1(n8986), .A2(n236), .Y(n8985) );
  AND2X1_RVT U8970 ( .A1(n8987), .A2(n8988), .Y(n8986) );
  OR2X1_RVT U8971 ( .A1(n12297), .A2(n8990), .Y(n8988) );
  OR2X1_RVT U8972 ( .A1(n8976), .A2(n8991), .Y(n8987) );
  OR2X1_RVT U8973 ( .A1(n8992), .A2(n12303), .Y(n8984) );
  AND2X1_RVT U8974 ( .A1(n8994), .A2(n8995), .Y(n8992) );
  OR2X1_RVT U8975 ( .A1(n8996), .A2(n8997), .Y(n8978) );
  AND2X1_RVT U8976 ( .A1(n8998), .A2(n8999), .Y(n8996) );
  OR2X1_RVT U8977 ( .A1(n12298), .A2(n9000), .Y(n8999) );
  AND2X1_RVT U8978 ( .A1(n9001), .A2(n9002), .Y(n8998) );
  AND2X1_RVT U8979 ( .A1(n9003), .A2(n9004), .Y(n8977) );
  OR2X1_RVT U8980 ( .A1(n9005), .A2(n12280), .Y(n9004) );
  AND2X1_RVT U8981 ( .A1(n9007), .A2(n9008), .Y(n9005) );
  OR2X1_RVT U8982 ( .A1(n9009), .A2(n9010), .Y(n9008) );
  OR2X1_RVT U8983 ( .A1(n12289), .A2(n12284), .Y(n9010) );
  OR2X1_RVT U8984 ( .A1(n9013), .A2(n9014), .Y(n9003) );
  AND2X1_RVT U8985 ( .A1(n9015), .A2(n9016), .Y(n9013) );
  AND2X1_RVT U8986 ( .A1(n9017), .A2(n9018), .Y(n9015) );
  AND4X1_RVT U8987 ( .A1(n9019), .A2(n9020), .A3(n9021), .A4(n9022), .Y(n8961)
         );
  AND4X1_RVT U8988 ( .A1(n9023), .A2(n9024), .A3(n9025), .A4(n9026), .Y(n9022)
         );
  OR2X1_RVT U8989 ( .A1(n9027), .A2(n12309), .Y(n9026) );
  AND4X1_RVT U8990 ( .A1(n9029), .A2(n9030), .A3(n9031), .A4(n9032), .Y(n9027)
         );
  OR2X1_RVT U8991 ( .A1(n9033), .A2(n9000), .Y(n9032) );
  OR2X1_RVT U8992 ( .A1(n9034), .A2(n12295), .Y(n9031) );
  OR2X1_RVT U8993 ( .A1(n9036), .A2(n12286), .Y(n9025) );
  AND4X1_RVT U8994 ( .A1(n9037), .A2(n9038), .A3(n9039), .A4(n9040), .Y(n9036)
         );
  OR2X1_RVT U8995 ( .A1(n9041), .A2(n9042), .Y(n9040) );
  OR2X1_RVT U8996 ( .A1(n12303), .A2(n12298), .Y(n9042) );
  AND2X1_RVT U8997 ( .A1(n9043), .A2(n9044), .Y(n9039) );
  OR2X1_RVT U8998 ( .A1(n12754), .A2(n9045), .Y(n9038) );
  OR2X1_RVT U8999 ( .A1(n9046), .A2(n9047), .Y(n9037) );
  AND2X1_RVT U9000 ( .A1(n9048), .A2(n9049), .Y(n9046) );
  OR2X1_RVT U9001 ( .A1(n12303), .A2(n9050), .Y(n9049) );
  OR2X1_RVT U9002 ( .A1(n8983), .A2(n9051), .Y(n9024) );
  OR2X1_RVT U9003 ( .A1(n9050), .A2(n9052), .Y(n9023) );
  OR2X1_RVT U9004 ( .A1(n9053), .A2(n9054), .Y(n9021) );
  OR2X1_RVT U9005 ( .A1(n9055), .A2(n9048), .Y(n9020) );
  OR2X1_RVT U9006 ( .A1(n9056), .A2(n9057), .Y(n9019) );
  AND4X1_RVT U9007 ( .A1(n9058), .A2(n9059), .A3(n9060), .A4(n9061), .Y(n8960)
         );
  AND2X1_RVT U9008 ( .A1(n9062), .A2(n9063), .Y(n9061) );
  OR2X1_RVT U9009 ( .A1(n9047), .A2(n9064), .Y(n9063) );
  AND2X1_RVT U9010 ( .A1(n9065), .A2(n9066), .Y(n9062) );
  OR2X1_RVT U9011 ( .A1(n9067), .A2(n8990), .Y(n9066) );
  OR2X1_RVT U9012 ( .A1(n8991), .A2(n9068), .Y(n9065) );
  OR2X1_RVT U9013 ( .A1(n234), .A2(n9069), .Y(n9060) );
  OR2X1_RVT U9014 ( .A1(n9070), .A2(n12293), .Y(n9059) );
  OR2X1_RVT U9015 ( .A1(n12296), .A2(n9072), .Y(n9058) );
  AND4X1_RVT U9016 ( .A1(n9074), .A2(n9075), .A3(n9076), .A4(n9077), .Y(n9073)
         );
  AND4X1_RVT U9017 ( .A1(n9078), .A2(n8969), .A3(n9079), .A4(n9080), .Y(n9077)
         );
  AND4X1_RVT U9018 ( .A1(n9081), .A2(n9082), .A3(n9083), .A4(n9084), .Y(n9080)
         );
  OR2X1_RVT U9019 ( .A1(n8990), .A2(n9085), .Y(n9084) );
  OR2X1_RVT U9020 ( .A1(n9086), .A2(n12308), .Y(n9085) );
  OR2X1_RVT U9021 ( .A1(n8991), .A2(n9087), .Y(n9083) );
  OR2X1_RVT U9022 ( .A1(n234), .A2(n12292), .Y(n9087) );
  OR2X1_RVT U9023 ( .A1(n9088), .A2(n9034), .Y(n9082) );
  AND2X1_RVT U9024 ( .A1(n9045), .A2(n9089), .Y(n9088) );
  OR2X1_RVT U9025 ( .A1(n9090), .A2(n9091), .Y(n9081) );
  AND2X1_RVT U9026 ( .A1(n9092), .A2(n9093), .Y(n9090) );
  AND2X1_RVT U9027 ( .A1(n9094), .A2(n9095), .Y(n9079) );
  OR2X1_RVT U9028 ( .A1(n9041), .A2(n9096), .Y(n9095) );
  OR2X1_RVT U9029 ( .A1(n9097), .A2(n12752), .Y(n9096) );
  OR2X1_RVT U9030 ( .A1(n9098), .A2(n9099), .Y(n9094) );
  OR2X1_RVT U9031 ( .A1(n9100), .A2(n12297), .Y(n9099) );
  OR2X1_RVT U9032 ( .A1(n8976), .A2(n9101), .Y(n8969) );
  AND4X1_RVT U9033 ( .A1(n9102), .A2(n9103), .A3(n9104), .A4(n9105), .Y(n9076)
         );
  AND4X1_RVT U9034 ( .A1(n9106), .A2(n9107), .A3(n9108), .A4(n9109), .Y(n9105)
         );
  OR2X1_RVT U9035 ( .A1(n9110), .A2(n12311), .Y(n9109) );
  AND2X1_RVT U9036 ( .A1(n9112), .A2(n9113), .Y(n9110) );
  OR2X1_RVT U9037 ( .A1(n12280), .A2(n8991), .Y(n9113) );
  OR2X1_RVT U9038 ( .A1(n9114), .A2(n8993), .Y(n9108) );
  AND2X1_RVT U9039 ( .A1(n9115), .A2(n9116), .Y(n9114) );
  OR2X1_RVT U9040 ( .A1(n9117), .A2(n12751), .Y(n9107) );
  AND2X1_RVT U9041 ( .A1(n9118), .A2(n9119), .Y(n9117) );
  OR2X1_RVT U9042 ( .A1(n9120), .A2(n9069), .Y(n9119) );
  AND2X1_RVT U9043 ( .A1(n12311), .A2(n12295), .Y(n9120) );
  OR2X1_RVT U9044 ( .A1(n9121), .A2(n12281), .Y(n9106) );
  AND2X1_RVT U9045 ( .A1(n9123), .A2(n9124), .Y(n9121) );
  OR2X1_RVT U9046 ( .A1(n9125), .A2(n12287), .Y(n9104) );
  AND2X1_RVT U9047 ( .A1(n9126), .A2(n9127), .Y(n9125) );
  OR2X1_RVT U9048 ( .A1(n12295), .A2(n9128), .Y(n9127) );
  AND2X1_RVT U9049 ( .A1(n9129), .A2(n9130), .Y(n9126) );
  OR2X1_RVT U9050 ( .A1(n9131), .A2(n9132), .Y(n9129) );
  OR2X1_RVT U9051 ( .A1(n8976), .A2(n9047), .Y(n9132) );
  OR2X1_RVT U9052 ( .A1(n9133), .A2(n12748), .Y(n9103) );
  AND2X1_RVT U9053 ( .A1(n9134), .A2(n9135), .Y(n9133) );
  OR2X1_RVT U9054 ( .A1(n9136), .A2(n9137), .Y(n9102) );
  AND2X1_RVT U9055 ( .A1(n9138), .A2(n9139), .Y(n9136) );
  AND2X1_RVT U9056 ( .A1(n9140), .A2(n9141), .Y(n9138) );
  OR2X1_RVT U9057 ( .A1(n236), .A2(n9069), .Y(n9141) );
  OR2X1_RVT U9058 ( .A1(n12305), .A2(n9034), .Y(n9140) );
  AND4X1_RVT U9059 ( .A1(n9142), .A2(n9143), .A3(n9144), .A4(n9145), .Y(n9075)
         );
  AND4X1_RVT U9060 ( .A1(n9146), .A2(n9147), .A3(n9148), .A4(n9149), .Y(n9145)
         );
  OR2X1_RVT U9061 ( .A1(n9069), .A2(n9068), .Y(n9149) );
  OR2X1_RVT U9062 ( .A1(n9000), .A2(n9150), .Y(n9148) );
  OR2X1_RVT U9063 ( .A1(n9033), .A2(n9151), .Y(n9147) );
  OR2X1_RVT U9064 ( .A1(n8976), .A2(n9152), .Y(n9146) );
  AND2X1_RVT U9065 ( .A1(n9153), .A2(n9154), .Y(n9144) );
  OR2X1_RVT U9066 ( .A1(n12306), .A2(n9155), .Y(n9154) );
  OR2X1_RVT U9067 ( .A1(n12285), .A2(n9052), .Y(n9153) );
  OR2X1_RVT U9068 ( .A1(n9156), .A2(n9011), .Y(n9143) );
  AND4X1_RVT U9069 ( .A1(n9157), .A2(n9158), .A3(n9159), .A4(n9160), .Y(n9156)
         );
  OR2X1_RVT U9070 ( .A1(n9161), .A2(n8976), .Y(n9159) );
  OR2X1_RVT U9071 ( .A1(n12740), .A2(n9162), .Y(n9158) );
  OR2X1_RVT U9072 ( .A1(n9163), .A2(n12748), .Y(n9157) );
  AND2X1_RVT U9073 ( .A1(n9054), .A2(n9164), .Y(n9163) );
  OR2X1_RVT U9074 ( .A1(n9056), .A2(n9165), .Y(n9142) );
  AND4X1_RVT U9075 ( .A1(n9166), .A2(n9167), .A3(n9168), .A4(n9169), .Y(n9074)
         );
  AND4X1_RVT U9076 ( .A1(n9170), .A2(n9171), .A3(n9172), .A4(n9173), .Y(n9169)
         );
  OR2X1_RVT U9077 ( .A1(n12744), .A2(n9174), .Y(n9173) );
  OR2X1_RVT U9078 ( .A1(n12745), .A2(n9175), .Y(n9172) );
  OR2X1_RVT U9079 ( .A1(n12742), .A2(n9176), .Y(n9171) );
  OR2X1_RVT U9080 ( .A1(n12279), .A2(n9177), .Y(n9170) );
  OR2X1_RVT U9081 ( .A1(n9178), .A2(n12286), .Y(n9167) );
  AND4X1_RVT U9082 ( .A1(n9180), .A2(n9181), .A3(n9182), .A4(n9183), .Y(n9179)
         );
  AND4X1_RVT U9083 ( .A1(n9184), .A2(n9185), .A3(n9186), .A4(n9187), .Y(n9183)
         );
  AND4X1_RVT U9084 ( .A1(n9188), .A2(n8965), .A3(n9135), .A4(n9189), .Y(n9187)
         );
  OR2X1_RVT U9085 ( .A1(n9190), .A2(n12739), .Y(n8965) );
  AND2X1_RVT U9086 ( .A1(n9191), .A2(n9192), .Y(n9190) );
  OR2X1_RVT U9087 ( .A1(n9009), .A2(n9193), .Y(n9192) );
  OR2X1_RVT U9088 ( .A1(n9194), .A2(n9091), .Y(n9191) );
  OR2X1_RVT U9089 ( .A1(n9195), .A2(n9050), .Y(n9188) );
  AND2X1_RVT U9090 ( .A1(n9196), .A2(n9197), .Y(n9195) );
  OR2X1_RVT U9091 ( .A1(n12744), .A2(n9034), .Y(n9197) );
  OR2X1_RVT U9092 ( .A1(n9198), .A2(n8993), .Y(n9186) );
  AND2X1_RVT U9093 ( .A1(n9199), .A2(n9200), .Y(n9198) );
  OR2X1_RVT U9094 ( .A1(n9201), .A2(n12750), .Y(n9200) );
  AND2X1_RVT U9095 ( .A1(n9041), .A2(n9202), .Y(n9201) );
  OR2X1_RVT U9096 ( .A1(n9203), .A2(n12306), .Y(n9185) );
  AND2X1_RVT U9097 ( .A1(n9204), .A2(n9205), .Y(n9203) );
  OR2X1_RVT U9098 ( .A1(n9034), .A2(n9000), .Y(n9205) );
  OR2X1_RVT U9099 ( .A1(n9206), .A2(n12289), .Y(n9184) );
  AND2X1_RVT U9100 ( .A1(n9118), .A2(n9207), .Y(n9206) );
  OR2X1_RVT U9101 ( .A1(n9047), .A2(n9208), .Y(n9118) );
  AND4X1_RVT U9102 ( .A1(n9209), .A2(n9210), .A3(n9211), .A4(n9212), .Y(n9182)
         );
  OR2X1_RVT U9103 ( .A1(n9213), .A2(n12296), .Y(n9212) );
  AND2X1_RVT U9104 ( .A1(n9214), .A2(n9215), .Y(n9213) );
  OR2X1_RVT U9105 ( .A1(n9091), .A2(n8991), .Y(n9215) );
  AND2X1_RVT U9106 ( .A1(n9216), .A2(n9217), .Y(n9214) );
  OR2X1_RVT U9107 ( .A1(n9131), .A2(n9193), .Y(n9216) );
  AND2X1_RVT U9108 ( .A1(n9218), .A2(n9219), .Y(n9211) );
  OR2X1_RVT U9109 ( .A1(n9220), .A2(n9122), .Y(n9219) );
  AND2X1_RVT U9110 ( .A1(n9221), .A2(n9030), .Y(n9220) );
  OR2X1_RVT U9111 ( .A1(n8976), .A2(n9091), .Y(n9030) );
  OR2X1_RVT U9112 ( .A1(n9222), .A2(n236), .Y(n9218) );
  AND2X1_RVT U9113 ( .A1(n9223), .A2(n9224), .Y(n9222) );
  OR2X1_RVT U9114 ( .A1(n9225), .A2(n12298), .Y(n9224) );
  AND2X1_RVT U9115 ( .A1(n9226), .A2(n9227), .Y(n9225) );
  OR2X1_RVT U9116 ( .A1(n12293), .A2(n9041), .Y(n9227) );
  OR2X1_RVT U9117 ( .A1(n12754), .A2(n12295), .Y(n9226) );
  AND2X1_RVT U9118 ( .A1(n9092), .A2(n9202), .Y(n9223) );
  OR2X1_RVT U9119 ( .A1(n9122), .A2(n9228), .Y(n9092) );
  OR2X1_RVT U9120 ( .A1(n12749), .A2(n12745), .Y(n9228) );
  OR2X1_RVT U9121 ( .A1(n9229), .A2(n9111), .Y(n9210) );
  AND4X1_RVT U9122 ( .A1(n9070), .A2(n9230), .A3(n9231), .A4(n9232), .Y(n9229)
         );
  OR2X1_RVT U9123 ( .A1(n12297), .A2(n9091), .Y(n9232) );
  AND2X1_RVT U9124 ( .A1(n9233), .A2(n9234), .Y(n9231) );
  OR2X1_RVT U9125 ( .A1(n12754), .A2(n12306), .Y(n9230) );
  AND2X1_RVT U9126 ( .A1(n9235), .A2(n9236), .Y(n9070) );
  OR2X1_RVT U9127 ( .A1(n9237), .A2(n234), .Y(n9236) );
  OR2X1_RVT U9128 ( .A1(n9034), .A2(n12739), .Y(n9235) );
  AND2X1_RVT U9129 ( .A1(n9238), .A2(n9239), .Y(n9209) );
  OR2X1_RVT U9130 ( .A1(n9240), .A2(n12741), .Y(n9239) );
  AND2X1_RVT U9131 ( .A1(n9241), .A2(n9242), .Y(n9240) );
  OR2X1_RVT U9132 ( .A1(n9243), .A2(n12300), .Y(n9242) );
  AND2X1_RVT U9133 ( .A1(n9244), .A2(n9245), .Y(n9243) );
  AND2X1_RVT U9134 ( .A1(n9246), .A2(n9247), .Y(n9241) );
  OR2X1_RVT U9135 ( .A1(n9248), .A2(n12309), .Y(n9238) );
  AND4X1_RVT U9136 ( .A1(n9249), .A2(n9250), .A3(n9251), .A4(n9252), .Y(n9248)
         );
  OR2X1_RVT U9137 ( .A1(n12753), .A2(n9253), .Y(n9251) );
  OR2X1_RVT U9138 ( .A1(n234), .A2(n9048), .Y(n9250) );
  OR2X1_RVT U9139 ( .A1(n9137), .A2(n9091), .Y(n9249) );
  AND4X1_RVT U9140 ( .A1(n9254), .A2(n9255), .A3(n9256), .A4(n9257), .Y(n9181)
         );
  AND2X1_RVT U9141 ( .A1(n9258), .A2(n9101), .Y(n9257) );
  OR2X1_RVT U9142 ( .A1(n12284), .A2(n9067), .Y(n9101) );
  AND2X1_RVT U9143 ( .A1(n9259), .A2(n9260), .Y(n9258) );
  OR2X1_RVT U9144 ( .A1(n9261), .A2(n9016), .Y(n9260) );
  OR2X1_RVT U9145 ( .A1(n9068), .A2(n9128), .Y(n9259) );
  OR2X1_RVT U9146 ( .A1(n234), .A2(n9262), .Y(n9256) );
  OR2X1_RVT U9147 ( .A1(n12752), .A2(n9263), .Y(n9255) );
  OR2X1_RVT U9148 ( .A1(n9137), .A2(n9264), .Y(n9254) );
  AND4X1_RVT U9149 ( .A1(n9265), .A2(n9266), .A3(n9267), .A4(n9268), .Y(n9180)
         );
  AND2X1_RVT U9150 ( .A1(n9269), .A2(n9270), .Y(n9268) );
  OR2X1_RVT U9151 ( .A1(n12279), .A2(n9271), .Y(n9270) );
  AND2X1_RVT U9152 ( .A1(n9272), .A2(n9273), .Y(n9269) );
  OR2X1_RVT U9153 ( .A1(n9033), .A2(n9043), .Y(n9273) );
  OR2X1_RVT U9154 ( .A1(n12300), .A2(n9093), .Y(n9043) );
  OR2X1_RVT U9155 ( .A1(n12286), .A2(n9274), .Y(n9272) );
  OR2X1_RVT U9156 ( .A1(n9014), .A2(n9007), .Y(n9267) );
  OR2X1_RVT U9157 ( .A1(n9100), .A2(n9275), .Y(n9007) );
  OR2X1_RVT U9158 ( .A1(n12748), .A2(n9276), .Y(n9266) );
  OR2X1_RVT U9159 ( .A1(n12298), .A2(n9134), .Y(n9265) );
  OR2X1_RVT U9160 ( .A1(n12739), .A2(n9196), .Y(n9134) );
  AND4X1_RVT U9161 ( .A1(n9278), .A2(n9279), .A3(n9280), .A4(n9281), .Y(n9277)
         );
  AND4X1_RVT U9162 ( .A1(n9282), .A2(n9283), .A3(n9284), .A4(n9285), .Y(n9281)
         );
  OR2X1_RVT U9163 ( .A1(n244), .A2(n9286), .Y(n9285) );
  OR2X1_RVT U9164 ( .A1(n9287), .A2(n12311), .Y(n9286) );
  AND2X1_RVT U9165 ( .A1(n12300), .A2(n9053), .Y(n9287) );
  AND2X1_RVT U9166 ( .A1(n8968), .A2(n9288), .Y(n9284) );
  OR2X1_RVT U9167 ( .A1(n12289), .A2(n9289), .Y(n8968) );
  OR2X1_RVT U9168 ( .A1(n244), .A2(n9047), .Y(n9289) );
  OR2X1_RVT U9169 ( .A1(n9290), .A2(n8976), .Y(n9283) );
  AND2X1_RVT U9170 ( .A1(n9291), .A2(n9292), .Y(n9290) );
  AND2X1_RVT U9171 ( .A1(n9293), .A2(n9294), .Y(n9282) );
  OR2X1_RVT U9172 ( .A1(n9295), .A2(n9296), .Y(n9294) );
  AND2X1_RVT U9173 ( .A1(n9297), .A2(n9057), .Y(n9295) );
  OR2X1_RVT U9174 ( .A1(n9298), .A2(n9048), .Y(n9293) );
  AND2X1_RVT U9175 ( .A1(n9233), .A2(n9067), .Y(n9298) );
  OR2X1_RVT U9176 ( .A1(n12287), .A2(n9299), .Y(n9233) );
  OR2X1_RVT U9177 ( .A1(n12754), .A2(n12297), .Y(n9299) );
  AND4X1_RVT U9178 ( .A1(n9300), .A2(n9301), .A3(n9302), .A4(n9303), .Y(n9280)
         );
  OR2X1_RVT U9179 ( .A1(n9304), .A2(n12744), .Y(n9303) );
  AND2X1_RVT U9180 ( .A1(n9116), .A2(n9305), .Y(n9304) );
  OR2X1_RVT U9181 ( .A1(n12752), .A2(n9161), .Y(n9116) );
  AND2X1_RVT U9182 ( .A1(n9306), .A2(n9307), .Y(n9302) );
  OR2X1_RVT U9183 ( .A1(n9308), .A2(n12742), .Y(n9307) );
  AND2X1_RVT U9184 ( .A1(n9309), .A2(n9310), .Y(n9308) );
  OR2X1_RVT U9185 ( .A1(n9011), .A2(n9253), .Y(n9310) );
  OR2X1_RVT U9186 ( .A1(n9311), .A2(n12740), .Y(n9306) );
  AND2X1_RVT U9187 ( .A1(n9312), .A2(n9313), .Y(n9311) );
  OR2X1_RVT U9188 ( .A1(n9314), .A2(n12300), .Y(n9301) );
  AND2X1_RVT U9189 ( .A1(n9315), .A2(n9316), .Y(n9314) );
  AND2X1_RVT U9190 ( .A1(n9317), .A2(n9318), .Y(n9315) );
  AND2X1_RVT U9191 ( .A1(n9319), .A2(n9320), .Y(n9300) );
  OR2X1_RVT U9192 ( .A1(n9321), .A2(n9237), .Y(n9320) );
  AND2X1_RVT U9193 ( .A1(n9322), .A2(n9068), .Y(n9321) );
  AND2X1_RVT U9194 ( .A1(n9323), .A2(n9324), .Y(n9322) );
  OR2X1_RVT U9195 ( .A1(n9325), .A2(n12303), .Y(n9319) );
  AND2X1_RVT U9196 ( .A1(n9326), .A2(n9327), .Y(n9325) );
  OR2X1_RVT U9197 ( .A1(n12751), .A2(n12305), .Y(n9327) );
  AND2X1_RVT U9198 ( .A1(n9057), .A2(n9328), .Y(n9326) );
  AND4X1_RVT U9199 ( .A1(n9329), .A2(n9330), .A3(n9331), .A4(n9332), .Y(n9279)
         );
  AND2X1_RVT U9200 ( .A1(n9333), .A2(n9334), .Y(n9332) );
  OR2X1_RVT U9201 ( .A1(n9050), .A2(n9124), .Y(n9334) );
  OR2X1_RVT U9202 ( .A1(n12746), .A2(n9057), .Y(n9124) );
  AND2X1_RVT U9203 ( .A1(n9335), .A2(n9336), .Y(n9333) );
  OR2X1_RVT U9204 ( .A1(n9202), .A2(n9016), .Y(n9336) );
  OR2X1_RVT U9205 ( .A1(n12753), .A2(n12296), .Y(n9016) );
  OR2X1_RVT U9206 ( .A1(n9100), .A2(n9150), .Y(n9335) );
  OR2X1_RVT U9207 ( .A1(n12741), .A2(n9337), .Y(n9150) );
  OR2X1_RVT U9208 ( .A1(n9338), .A2(n12279), .Y(n9331) );
  AND4X1_RVT U9209 ( .A1(n9339), .A2(n9340), .A3(n9341), .A4(n9342), .Y(n9338)
         );
  OR2X1_RVT U9210 ( .A1(n9275), .A2(n9048), .Y(n9341) );
  OR2X1_RVT U9211 ( .A1(n9343), .A2(n9045), .Y(n9340) );
  OR2X1_RVT U9212 ( .A1(n12750), .A2(n9000), .Y(n9339) );
  OR2X1_RVT U9213 ( .A1(n9344), .A2(n12280), .Y(n9330) );
  AND2X1_RVT U9214 ( .A1(n9345), .A2(n9346), .Y(n9344) );
  OR2X1_RVT U9215 ( .A1(n9275), .A2(n9000), .Y(n9346) );
  AND2X1_RVT U9216 ( .A1(n9347), .A2(n9276), .Y(n9345) );
  OR2X1_RVT U9217 ( .A1(n9048), .A2(n9348), .Y(n9276) );
  OR2X1_RVT U9218 ( .A1(n12741), .A2(n12753), .Y(n9348) );
  OR2X1_RVT U9219 ( .A1(n9349), .A2(n12287), .Y(n9329) );
  AND4X1_RVT U9220 ( .A1(n9350), .A2(n9263), .A3(n9072), .A4(n9044), .Y(n9349)
         );
  OR2X1_RVT U9221 ( .A1(n9069), .A2(n9351), .Y(n9044) );
  OR2X1_RVT U9222 ( .A1(n12743), .A2(n9006), .Y(n9351) );
  OR2X1_RVT U9223 ( .A1(n9131), .A2(n9165), .Y(n9072) );
  OR2X1_RVT U9224 ( .A1(n9050), .A2(n9352), .Y(n9263) );
  OR2X1_RVT U9225 ( .A1(n12311), .A2(n12280), .Y(n9352) );
  OR2X1_RVT U9226 ( .A1(n9009), .A2(n9353), .Y(n9350) );
  OR2X1_RVT U9227 ( .A1(n9354), .A2(n12285), .Y(n9353) );
  AND4X1_RVT U9228 ( .A1(n9355), .A2(n9356), .A3(n9357), .A4(n9358), .Y(n9278)
         );
  AND2X1_RVT U9229 ( .A1(n9359), .A2(n9360), .Y(n9358) );
  AND2X1_RVT U9230 ( .A1(n9361), .A2(n9362), .Y(n9359) );
  OR2X1_RVT U9231 ( .A1(n9041), .A2(n9316), .Y(n9362) );
  OR2X1_RVT U9232 ( .A1(n9053), .A2(n9363), .Y(n9316) );
  OR2X1_RVT U9233 ( .A1(n12742), .A2(n12744), .Y(n9363) );
  OR2X1_RVT U9234 ( .A1(n12749), .A2(n9364), .Y(n9361) );
  OR2X1_RVT U9235 ( .A1(n12296), .A2(n9365), .Y(n9357) );
  OR2X1_RVT U9236 ( .A1(n12752), .A2(n9366), .Y(n9356) );
  OR2X1_RVT U9237 ( .A1(n9053), .A2(n9367), .Y(n9355) );
  AND4X1_RVT U9238 ( .A1(n9369), .A2(n9370), .A3(n9371), .A4(n9372), .Y(n9368)
         );
  AND4X1_RVT U9239 ( .A1(n9373), .A2(n9374), .A3(n9375), .A4(n9376), .Y(n9372)
         );
  AND4X1_RVT U9240 ( .A1(n9377), .A2(n9378), .A3(n8970), .A4(n9379), .Y(n9376)
         );
  OR2X1_RVT U9241 ( .A1(n9111), .A2(n9380), .Y(n8970) );
  OR2X1_RVT U9242 ( .A1(n9202), .A2(n236), .Y(n9380) );
  OR2X1_RVT U9243 ( .A1(n8974), .A2(n9381), .Y(n9378) );
  OR2X1_RVT U9244 ( .A1(n12747), .A2(n12750), .Y(n9381) );
  OR2X1_RVT U9245 ( .A1(n9237), .A2(n9382), .Y(n9377) );
  OR2X1_RVT U9246 ( .A1(n9383), .A2(n9011), .Y(n9382) );
  AND2X1_RVT U9247 ( .A1(n12300), .A2(n9111), .Y(n9383) );
  OR2X1_RVT U9248 ( .A1(n9384), .A2(n12306), .Y(n9375) );
  AND2X1_RVT U9249 ( .A1(n9252), .A2(n9324), .Y(n9384) );
  OR2X1_RVT U9250 ( .A1(n236), .A2(n9385), .Y(n9324) );
  OR2X1_RVT U9251 ( .A1(n12279), .A2(n12746), .Y(n9385) );
  OR2X1_RVT U9252 ( .A1(n9041), .A2(n9386), .Y(n9252) );
  OR2X1_RVT U9253 ( .A1(n12744), .A2(n9033), .Y(n9386) );
  OR2X1_RVT U9254 ( .A1(n9387), .A2(n8991), .Y(n9374) );
  AND2X1_RVT U9255 ( .A1(n9388), .A2(n9196), .Y(n9387) );
  OR2X1_RVT U9256 ( .A1(n9097), .A2(n9091), .Y(n9373) );
  AND4X1_RVT U9257 ( .A1(n9389), .A2(n9390), .A3(n9391), .A4(n9392), .Y(n9371)
         );
  AND2X1_RVT U9258 ( .A1(n9393), .A2(n9394), .Y(n9392) );
  OR2X1_RVT U9259 ( .A1(n9395), .A2(n12300), .Y(n9394) );
  AND2X1_RVT U9260 ( .A1(n9396), .A2(n9064), .Y(n9395) );
  AND2X1_RVT U9261 ( .A1(n9397), .A2(n9398), .Y(n9393) );
  OR2X1_RVT U9262 ( .A1(n9399), .A2(n9047), .Y(n9398) );
  AND2X1_RVT U9263 ( .A1(n9018), .A2(n8990), .Y(n9399) );
  OR2X1_RVT U9264 ( .A1(n12752), .A2(n9089), .Y(n9018) );
  OR2X1_RVT U9265 ( .A1(n9400), .A2(n9100), .Y(n9397) );
  AND2X1_RVT U9266 ( .A1(n9292), .A2(n9401), .Y(n9400) );
  OR2X1_RVT U9267 ( .A1(n12753), .A2(n9128), .Y(n9292) );
  OR2X1_RVT U9268 ( .A1(n9402), .A2(n12744), .Y(n9391) );
  AND2X1_RVT U9269 ( .A1(n8995), .A2(n9403), .Y(n9402) );
  OR2X1_RVT U9270 ( .A1(n9131), .A2(n9055), .Y(n9403) );
  OR2X1_RVT U9271 ( .A1(n9034), .A2(n9237), .Y(n8995) );
  OR2X1_RVT U9272 ( .A1(n9404), .A2(n234), .Y(n9390) );
  AND2X1_RVT U9273 ( .A1(n9045), .A2(n9405), .Y(n9404) );
  OR2X1_RVT U9274 ( .A1(n9406), .A2(n12284), .Y(n9405) );
  AND2X1_RVT U9275 ( .A1(n9407), .A2(n9408), .Y(n9406) );
  OR2X1_RVT U9276 ( .A1(n12745), .A2(n9028), .Y(n9408) );
  OR2X1_RVT U9277 ( .A1(n12311), .A2(n9131), .Y(n9045) );
  OR2X1_RVT U9278 ( .A1(n9409), .A2(n9115), .Y(n9389) );
  AND2X1_RVT U9279 ( .A1(n9048), .A2(n9093), .Y(n9409) );
  OR2X1_RVT U9280 ( .A1(n12741), .A2(n8976), .Y(n9093) );
  AND4X1_RVT U9281 ( .A1(n9410), .A2(n9411), .A3(n9412), .A4(n9413), .Y(n9370)
         );
  AND4X1_RVT U9282 ( .A1(n9414), .A2(n9415), .A3(n9416), .A4(n9417), .Y(n9413)
         );
  OR2X1_RVT U9283 ( .A1(n9418), .A2(n12752), .Y(n9417) );
  AND2X1_RVT U9284 ( .A1(n9151), .A2(n9419), .Y(n9418) );
  OR2X1_RVT U9285 ( .A1(n12308), .A2(n9000), .Y(n9419) );
  OR2X1_RVT U9286 ( .A1(n9420), .A2(n8993), .Y(n9416) );
  AND2X1_RVT U9287 ( .A1(n9421), .A2(n9422), .Y(n9420) );
  OR2X1_RVT U9288 ( .A1(n9423), .A2(n9028), .Y(n9422) );
  AND2X1_RVT U9289 ( .A1(n9053), .A2(n9041), .Y(n9423) );
  AND2X1_RVT U9290 ( .A1(n9055), .A2(n9297), .Y(n9421) );
  OR2X1_RVT U9291 ( .A1(n12309), .A2(n9193), .Y(n9297) );
  OR2X1_RVT U9292 ( .A1(n9424), .A2(n12298), .Y(n9415) );
  AND2X1_RVT U9293 ( .A1(n9425), .A2(n9426), .Y(n9424) );
  OR2X1_RVT U9294 ( .A1(n9041), .A2(n9427), .Y(n9426) );
  AND2X1_RVT U9295 ( .A1(n9123), .A2(n9317), .Y(n9425) );
  OR2X1_RVT U9296 ( .A1(n9033), .A2(n9208), .Y(n9317) );
  OR2X1_RVT U9297 ( .A1(n9006), .A2(n9428), .Y(n9123) );
  OR2X1_RVT U9298 ( .A1(n9429), .A2(n8976), .Y(n9414) );
  AND4X1_RVT U9299 ( .A1(n9430), .A2(n9431), .A3(n9432), .A4(n9365), .Y(n9429)
         );
  OR2X1_RVT U9300 ( .A1(n9069), .A2(n9433), .Y(n9365) );
  OR2X1_RVT U9301 ( .A1(n12279), .A2(n9033), .Y(n9433) );
  OR2X1_RVT U9302 ( .A1(n12749), .A2(n9275), .Y(n9431) );
  OR2X1_RVT U9303 ( .A1(n9034), .A2(n9131), .Y(n9430) );
  OR2X1_RVT U9304 ( .A1(n9202), .A2(n9244), .Y(n9412) );
  OR2X1_RVT U9305 ( .A1(n9434), .A2(n12282), .Y(n9411) );
  AND4X1_RVT U9306 ( .A1(n9435), .A2(n9436), .A3(n9078), .A4(n9176), .Y(n9434)
         );
  OR2X1_RVT U9307 ( .A1(n9000), .A2(n9165), .Y(n9176) );
  OR2X1_RVT U9308 ( .A1(n12749), .A2(n234), .Y(n9165) );
  OR2X1_RVT U9309 ( .A1(n8993), .A2(n9057), .Y(n9078) );
  OR2X1_RVT U9310 ( .A1(n12741), .A2(n9428), .Y(n9410) );
  AND4X1_RVT U9311 ( .A1(n9437), .A2(n9438), .A3(n9439), .A4(n9440), .Y(n9369)
         );
  OR2X1_RVT U9312 ( .A1(n12287), .A2(n9441), .Y(n9440) );
  AND2X1_RVT U9313 ( .A1(n9442), .A2(n9443), .Y(n9439) );
  OR2X1_RVT U9314 ( .A1(n12308), .A2(n9196), .Y(n9443) );
  OR2X1_RVT U9315 ( .A1(n8983), .A2(n9057), .Y(n9442) );
  OR2X1_RVT U9316 ( .A1(n236), .A2(n9014), .Y(n9057) );
  OR2X1_RVT U9317 ( .A1(n12311), .A2(n9175), .Y(n9438) );
  OR2X1_RVT U9318 ( .A1(n9050), .A2(n9444), .Y(n9175) );
  AND2X1_RVT U9319 ( .A1(n9445), .A2(n9446), .Y(n9437) );
  OR2X1_RVT U9320 ( .A1(n12280), .A2(n9447), .Y(n9446) );
  OR2X1_RVT U9321 ( .A1(n9053), .A2(n9002), .Y(n9445) );
  OR2X1_RVT U9322 ( .A1(n8976), .A2(n9261), .Y(n9002) );
  AND4X1_RVT U9323 ( .A1(n9449), .A2(n9450), .A3(n9451), .A4(n9452), .Y(n9448)
         );
  AND4X1_RVT U9324 ( .A1(n9453), .A2(n9454), .A3(n9455), .A4(n9456), .Y(n9452)
         );
  AND4X1_RVT U9325 ( .A1(n9189), .A2(n9379), .A3(n9457), .A4(n9458), .Y(n9456)
         );
  OR2X1_RVT U9326 ( .A1(n9459), .A2(n9460), .Y(n9379) );
  OR2X1_RVT U9327 ( .A1(n8974), .A2(n9244), .Y(n9189) );
  OR2X1_RVT U9328 ( .A1(n12750), .A2(n12296), .Y(n9244) );
  AND4X1_RVT U9329 ( .A1(n9447), .A2(n9313), .A3(n9436), .A4(n8971), .Y(n9455)
         );
  OR2X1_RVT U9330 ( .A1(n9461), .A2(n9161), .Y(n8971) );
  OR2X1_RVT U9331 ( .A1(n8976), .A2(n9462), .Y(n9436) );
  OR2X1_RVT U9332 ( .A1(n9009), .A2(n234), .Y(n9313) );
  OR2X1_RVT U9333 ( .A1(n9000), .A2(n9463), .Y(n9447) );
  OR2X1_RVT U9334 ( .A1(n12286), .A2(n12306), .Y(n9463) );
  AND4X1_RVT U9335 ( .A1(n9464), .A2(n9465), .A3(n9466), .A4(n9467), .Y(n9454)
         );
  OR2X1_RVT U9336 ( .A1(n9253), .A2(n9468), .Y(n9467) );
  OR2X1_RVT U9337 ( .A1(n12306), .A2(n9033), .Y(n9468) );
  OR2X1_RVT U9338 ( .A1(n9162), .A2(n9469), .Y(n9466) );
  OR2X1_RVT U9339 ( .A1(n12751), .A2(n9050), .Y(n9469) );
  OR2X1_RVT U9340 ( .A1(n9388), .A2(n9470), .Y(n9465) );
  OR2X1_RVT U9341 ( .A1(n9471), .A2(n9047), .Y(n9470) );
  OR2X1_RVT U9342 ( .A1(n12303), .A2(n9472), .Y(n9464) );
  OR2X1_RVT U9343 ( .A1(n9473), .A2(n12286), .Y(n9472) );
  AND2X1_RVT U9344 ( .A1(n9261), .A2(n9474), .Y(n9473) );
  AND2X1_RVT U9345 ( .A1(n9475), .A2(n9476), .Y(n9453) );
  OR2X1_RVT U9346 ( .A1(n9477), .A2(n9028), .Y(n9476) );
  AND2X1_RVT U9347 ( .A1(n9478), .A2(n9479), .Y(n9477) );
  OR2X1_RVT U9348 ( .A1(n12285), .A2(n9221), .Y(n9479) );
  OR2X1_RVT U9349 ( .A1(n12289), .A2(n9296), .Y(n9478) );
  AND2X1_RVT U9350 ( .A1(n9480), .A2(n9481), .Y(n9475) );
  OR2X1_RVT U9351 ( .A1(n9482), .A2(n9067), .Y(n9481) );
  AND2X1_RVT U9352 ( .A1(n9483), .A2(n9484), .Y(n9482) );
  OR2X1_RVT U9353 ( .A1(n12292), .A2(n244), .Y(n9484) );
  NAND2X1_RVT U9354 ( .A1(n9050), .A2(n12743), .Y(n9483) );
  OR2X1_RVT U9355 ( .A1(n9485), .A2(n236), .Y(n9480) );
  AND2X1_RVT U9356 ( .A1(n9274), .A2(n9151), .Y(n9485) );
  OR2X1_RVT U9357 ( .A1(n9000), .A2(n9486), .Y(n9151) );
  OR2X1_RVT U9358 ( .A1(n12754), .A2(n12281), .Y(n9486) );
  AND4X1_RVT U9359 ( .A1(n9168), .A2(n9487), .A3(n9360), .A4(n9488), .Y(n9451)
         );
  AND4X1_RVT U9360 ( .A1(n9489), .A2(n9490), .A3(n9491), .A4(n9492), .Y(n9488)
         );
  OR2X1_RVT U9361 ( .A1(n9131), .A2(n9052), .Y(n9492) );
  OR2X1_RVT U9362 ( .A1(n9069), .A2(n9098), .Y(n9491) );
  OR2X1_RVT U9363 ( .A1(n12742), .A2(n9323), .Y(n9490) );
  OR2X1_RVT U9364 ( .A1(n9047), .A2(n9029), .Y(n9323) );
  OR2X1_RVT U9365 ( .A1(n12750), .A2(n9111), .Y(n9029) );
  OR2X1_RVT U9366 ( .A1(n12295), .A2(n9152), .Y(n9489) );
  OR2X1_RVT U9367 ( .A1(n9033), .A2(n9261), .Y(n9152) );
  OR2X1_RVT U9368 ( .A1(n12279), .A2(n9237), .Y(n9261) );
  AND2X1_RVT U9369 ( .A1(n9493), .A2(n9494), .Y(n9360) );
  OR2X1_RVT U9370 ( .A1(n9495), .A2(n9100), .Y(n9494) );
  OR2X1_RVT U9371 ( .A1(n12305), .A2(n236), .Y(n9495) );
  OR2X1_RVT U9372 ( .A1(n9496), .A2(n8983), .Y(n9493) );
  OR2X1_RVT U9373 ( .A1(n12741), .A2(n9100), .Y(n8983) );
  OR2X1_RVT U9374 ( .A1(n8997), .A2(n9047), .Y(n9496) );
  OR2X1_RVT U9375 ( .A1(n12287), .A2(n9366), .Y(n9487) );
  AND2X1_RVT U9376 ( .A1(n9497), .A2(n9498), .Y(n9168) );
  OR2X1_RVT U9377 ( .A1(n9051), .A2(n9089), .Y(n9498) );
  OR2X1_RVT U9378 ( .A1(n9499), .A2(n9500), .Y(n9497) );
  AND4X1_RVT U9379 ( .A1(n9501), .A2(n9502), .A3(n9503), .A4(n9504), .Y(n9450)
         );
  OR2X1_RVT U9380 ( .A1(n9505), .A2(n9237), .Y(n9504) );
  AND2X1_RVT U9381 ( .A1(n9506), .A2(n9246), .Y(n9505) );
  OR2X1_RVT U9382 ( .A1(n12293), .A2(n9462), .Y(n9246) );
  OR2X1_RVT U9383 ( .A1(n9507), .A2(n12747), .Y(n9503) );
  AND2X1_RVT U9384 ( .A1(n9174), .A2(n9139), .Y(n9507) );
  OR2X1_RVT U9385 ( .A1(n12741), .A2(n9115), .Y(n9139) );
  OR2X1_RVT U9386 ( .A1(n9508), .A2(n9194), .Y(n9502) );
  AND2X1_RVT U9387 ( .A1(n9509), .A2(n9510), .Y(n9508) );
  OR2X1_RVT U9388 ( .A1(n12282), .A2(n9053), .Y(n9510) );
  AND2X1_RVT U9389 ( .A1(n9511), .A2(n9091), .Y(n9509) );
  OR2X1_RVT U9390 ( .A1(n234), .A2(n9050), .Y(n9511) );
  OR2X1_RVT U9391 ( .A1(n9512), .A2(n8991), .Y(n9501) );
  AND2X1_RVT U9392 ( .A1(n9513), .A2(n9514), .Y(n9512) );
  NAND2X1_RVT U9393 ( .A1(n8976), .A2(n9354), .Y(n9514) );
  AND2X1_RVT U9394 ( .A1(n9515), .A2(n9204), .Y(n9513) );
  OR2X1_RVT U9395 ( .A1(n9137), .A2(n9462), .Y(n9204) );
  OR2X1_RVT U9396 ( .A1(n12302), .A2(n9516), .Y(n9515) );
  AND4X1_RVT U9397 ( .A1(n9517), .A2(n9518), .A3(n9519), .A4(n9520), .Y(n9449)
         );
  OR2X1_RVT U9398 ( .A1(n9521), .A2(n9014), .Y(n9520) );
  AND2X1_RVT U9399 ( .A1(n9522), .A2(n9155), .Y(n9521) );
  AND2X1_RVT U9400 ( .A1(n9523), .A2(n9177), .Y(n9522) );
  OR2X1_RVT U9401 ( .A1(n236), .A2(n9500), .Y(n9177) );
  OR2X1_RVT U9402 ( .A1(n12281), .A2(n9111), .Y(n9500) );
  OR2X1_RVT U9403 ( .A1(n9524), .A2(n12298), .Y(n9519) );
  AND2X1_RVT U9404 ( .A1(n9525), .A2(n9526), .Y(n9524) );
  OR2X1_RVT U9405 ( .A1(n9527), .A2(n12739), .Y(n9526) );
  AND2X1_RVT U9406 ( .A1(n9528), .A2(n9529), .Y(n9527) );
  OR2X1_RVT U9407 ( .A1(n12280), .A2(n9388), .Y(n9529) );
  OR2X1_RVT U9408 ( .A1(n12746), .A2(n9034), .Y(n9528) );
  AND2X1_RVT U9409 ( .A1(n9530), .A2(n9531), .Y(n9525) );
  OR2X1_RVT U9410 ( .A1(n9000), .A2(n9532), .Y(n9530) );
  OR2X1_RVT U9411 ( .A1(n9533), .A2(n9034), .Y(n9518) );
  AND4X1_RVT U9412 ( .A1(n9534), .A2(n9535), .A3(n9536), .A4(n9000), .Y(n9533)
         );
  OR2X1_RVT U9413 ( .A1(n12747), .A2(n9050), .Y(n9536) );
  OR2X1_RVT U9414 ( .A1(n12292), .A2(n9069), .Y(n9535) );
  OR2X1_RVT U9415 ( .A1(n9122), .A2(n9100), .Y(n9534) );
  OR2X1_RVT U9416 ( .A1(n9537), .A2(n8976), .Y(n9517) );
  AND4X1_RVT U9417 ( .A1(n9401), .A2(n9538), .A3(n9199), .A4(n9115), .Y(n9537)
         );
  OR2X1_RVT U9418 ( .A1(n9069), .A2(n9532), .Y(n9199) );
  OR2X1_RVT U9419 ( .A1(n9237), .A2(n9444), .Y(n9538) );
  OR2X1_RVT U9420 ( .A1(n12286), .A2(n9202), .Y(n9401) );
  AND4X1_RVT U9421 ( .A1(n9540), .A2(n9541), .A3(n9542), .A4(n9543), .Y(n9539)
         );
  AND4X1_RVT U9422 ( .A1(n9052), .A2(n9288), .A3(n9544), .A4(n9545), .Y(n9543)
         );
  AND4X1_RVT U9423 ( .A1(n9367), .A2(n9312), .A3(n9457), .A4(n9458), .Y(n9545)
         );
  OR2X1_RVT U9424 ( .A1(n9460), .A2(n8973), .Y(n9458) );
  OR2X1_RVT U9425 ( .A1(n12745), .A2(n9091), .Y(n8973) );
  OR2X1_RVT U9426 ( .A1(n8990), .A2(n9499), .Y(n9457) );
  OR2X1_RVT U9427 ( .A1(n12750), .A2(n12300), .Y(n9499) );
  OR2X1_RVT U9428 ( .A1(n12739), .A2(n9111), .Y(n8990) );
  OR2X1_RVT U9429 ( .A1(n12751), .A2(n9009), .Y(n9312) );
  OR2X1_RVT U9430 ( .A1(n12309), .A2(n12293), .Y(n9009) );
  OR2X1_RVT U9431 ( .A1(n9131), .A2(n9546), .Y(n9367) );
  OR2X1_RVT U9432 ( .A1(n12300), .A2(n9035), .Y(n9546) );
  OR2X1_RVT U9433 ( .A1(n9033), .A2(n9547), .Y(n9544) );
  OR2X1_RVT U9434 ( .A1(n9161), .A2(n12291), .Y(n9547) );
  OR2X1_RVT U9435 ( .A1(n9100), .A2(n9548), .Y(n9288) );
  OR2X1_RVT U9436 ( .A1(n9034), .A2(n12298), .Y(n9548) );
  OR2X1_RVT U9437 ( .A1(n12743), .A2(n9459), .Y(n9052) );
  OR2X1_RVT U9438 ( .A1(n12293), .A2(n9051), .Y(n9459) );
  AND4X1_RVT U9439 ( .A1(n9549), .A2(n9550), .A3(n9551), .A4(n9552), .Y(n9542)
         );
  AND4X1_RVT U9440 ( .A1(n9553), .A2(n9554), .A3(n9555), .A4(n9556), .Y(n9552)
         );
  OR2X1_RVT U9441 ( .A1(n9067), .A2(n9557), .Y(n9556) );
  OR2X1_RVT U9442 ( .A1(n12282), .A2(n9137), .Y(n9557) );
  OR2X1_RVT U9443 ( .A1(n9050), .A2(n9558), .Y(n9555) );
  OR2X1_RVT U9444 ( .A1(n9559), .A2(n9014), .Y(n9558) );
  AND2X1_RVT U9445 ( .A1(n8993), .A2(n9053), .Y(n9559) );
  OR2X1_RVT U9446 ( .A1(n9560), .A2(n9561), .Y(n9554) );
  AND2X1_RVT U9447 ( .A1(n9208), .A2(n9164), .Y(n9560) );
  OR2X1_RVT U9448 ( .A1(n12744), .A2(n244), .Y(n9164) );
  OR2X1_RVT U9449 ( .A1(n12740), .A2(n12303), .Y(n9208) );
  OR2X1_RVT U9450 ( .A1(n9562), .A2(n9048), .Y(n9553) );
  AND2X1_RVT U9451 ( .A1(n9444), .A2(n9563), .Y(n9562) );
  OR2X1_RVT U9452 ( .A1(n12742), .A2(n236), .Y(n9563) );
  OR2X1_RVT U9453 ( .A1(n9564), .A2(n12305), .Y(n9551) );
  AND2X1_RVT U9454 ( .A1(n9435), .A2(n9565), .Y(n9564) );
  OR2X1_RVT U9455 ( .A1(n9041), .A2(n9388), .Y(n9565) );
  OR2X1_RVT U9456 ( .A1(n12286), .A2(n9253), .Y(n9435) );
  OR2X1_RVT U9457 ( .A1(n12746), .A2(n9041), .Y(n9253) );
  OR2X1_RVT U9458 ( .A1(n9566), .A2(n9202), .Y(n9550) );
  AND2X1_RVT U9459 ( .A1(n9155), .A2(n9427), .Y(n9566) );
  OR2X1_RVT U9460 ( .A1(n9011), .A2(n9100), .Y(n9155) );
  OR2X1_RVT U9461 ( .A1(n9567), .A2(n9091), .Y(n9549) );
  AND2X1_RVT U9462 ( .A1(n9054), .A2(n9056), .Y(n9567) );
  AND4X1_RVT U9463 ( .A1(n9568), .A2(n9569), .A3(n9570), .A4(n9571), .Y(n9541)
         );
  AND4X1_RVT U9464 ( .A1(n9572), .A2(n9573), .A3(n9574), .A4(n9575), .Y(n9571)
         );
  OR2X1_RVT U9465 ( .A1(n9576), .A2(n12289), .Y(n9575) );
  AND2X1_RVT U9466 ( .A1(n8982), .A2(n9274), .Y(n9576) );
  OR2X1_RVT U9467 ( .A1(n9131), .A2(n9162), .Y(n9274) );
  OR2X1_RVT U9468 ( .A1(n12292), .A2(n9014), .Y(n9162) );
  OR2X1_RVT U9469 ( .A1(n12296), .A2(n9577), .Y(n8982) );
  OR2X1_RVT U9470 ( .A1(n12279), .A2(n12285), .Y(n9577) );
  OR2X1_RVT U9471 ( .A1(n9578), .A2(n12303), .Y(n9574) );
  AND2X1_RVT U9472 ( .A1(n9291), .A2(n9579), .Y(n9578) );
  OR2X1_RVT U9473 ( .A1(n12308), .A2(n234), .Y(n9579) );
  OR2X1_RVT U9474 ( .A1(n12306), .A2(n9098), .Y(n9291) );
  OR2X1_RVT U9475 ( .A1(n9580), .A2(n12284), .Y(n9573) );
  AND2X1_RVT U9476 ( .A1(n9309), .A2(n9581), .Y(n9580) );
  OR2X1_RVT U9477 ( .A1(n12309), .A2(n9034), .Y(n9581) );
  OR2X1_RVT U9478 ( .A1(n8976), .A2(n9582), .Y(n9309) );
  OR2X1_RVT U9479 ( .A1(n9583), .A2(n9035), .Y(n9572) );
  AND2X1_RVT U9480 ( .A1(n9584), .A2(n9585), .Y(n9583) );
  OR2X1_RVT U9481 ( .A1(n9091), .A2(n12306), .Y(n9585) );
  AND2X1_RVT U9482 ( .A1(n9586), .A2(n9067), .Y(n9584) );
  OR2X1_RVT U9483 ( .A1(n9053), .A2(n9014), .Y(n9067) );
  OR2X1_RVT U9484 ( .A1(n12281), .A2(n9098), .Y(n9586) );
  OR2X1_RVT U9485 ( .A1(n12754), .A2(n9053), .Y(n9098) );
  OR2X1_RVT U9486 ( .A1(n9587), .A2(n9111), .Y(n9570) );
  AND4X1_RVT U9487 ( .A1(n9588), .A2(n9589), .A3(n9264), .A4(n9174), .Y(n9587)
         );
  OR2X1_RVT U9488 ( .A1(n9237), .A2(n9337), .Y(n9174) );
  OR2X1_RVT U9489 ( .A1(n9069), .A2(n9516), .Y(n9264) );
  OR2X1_RVT U9490 ( .A1(n12287), .A2(n12280), .Y(n9516) );
  OR2X1_RVT U9491 ( .A1(n236), .A2(n8991), .Y(n9589) );
  OR2X1_RVT U9492 ( .A1(n234), .A2(n12306), .Y(n9588) );
  OR2X1_RVT U9493 ( .A1(n9590), .A2(n9047), .Y(n9569) );
  AND2X1_RVT U9494 ( .A1(n9591), .A2(n9068), .Y(n9590) );
  AND2X1_RVT U9495 ( .A1(n9523), .A2(n9318), .Y(n9591) );
  OR2X1_RVT U9496 ( .A1(n9592), .A2(n12751), .Y(n9318) );
  AND2X1_RVT U9497 ( .A1(n9089), .A2(n9593), .Y(n9592) );
  OR2X1_RVT U9498 ( .A1(n12284), .A2(n8976), .Y(n9593) );
  OR2X1_RVT U9499 ( .A1(n9137), .A2(n9275), .Y(n9523) );
  OR2X1_RVT U9500 ( .A1(n9122), .A2(n9011), .Y(n9275) );
  OR2X1_RVT U9501 ( .A1(n9594), .A2(n9115), .Y(n9568) );
  AND2X1_RVT U9502 ( .A1(n9595), .A2(n12292), .Y(n9594) );
  AND2X1_RVT U9503 ( .A1(n9596), .A2(n9296), .Y(n9595) );
  OR2X1_RVT U9504 ( .A1(n9137), .A2(n9237), .Y(n9596) );
  AND4X1_RVT U9505 ( .A1(n9597), .A2(n9598), .A3(n9599), .A4(n9600), .Y(n9540)
         );
  AND2X1_RVT U9506 ( .A1(n9601), .A2(n9602), .Y(n9600) );
  OR2X1_RVT U9507 ( .A1(n12747), .A2(n9217), .Y(n9602) );
  OR2X1_RVT U9508 ( .A1(n12300), .A2(n9603), .Y(n9217) );
  OR2X1_RVT U9509 ( .A1(n9033), .A2(n9122), .Y(n9603) );
  AND2X1_RVT U9510 ( .A1(n9604), .A2(n9605), .Y(n9601) );
  OR2X1_RVT U9511 ( .A1(n9006), .A2(n9017), .Y(n9605) );
  OR2X1_RVT U9512 ( .A1(n9050), .A2(n9245), .Y(n9017) );
  OR2X1_RVT U9513 ( .A1(n12743), .A2(n9011), .Y(n9245) );
  OR2X1_RVT U9514 ( .A1(n9053), .A2(n9130), .Y(n9604) );
  OR2X1_RVT U9515 ( .A1(n9041), .A2(n9606), .Y(n9130) );
  OR2X1_RVT U9516 ( .A1(n9041), .A2(n9221), .Y(n9599) );
  OR2X1_RVT U9517 ( .A1(n236), .A2(n12302), .Y(n9221) );
  OR2X1_RVT U9518 ( .A1(n9607), .A2(n8997), .Y(n9598) );
  AND4X1_RVT U9519 ( .A1(n9608), .A2(n9609), .A3(n9610), .A4(n9611), .Y(n9607)
         );
  OR2X1_RVT U9520 ( .A1(n12741), .A2(n9612), .Y(n9610) );
  OR2X1_RVT U9521 ( .A1(n9613), .A2(n12748), .Y(n9612) );
  AND2X1_RVT U9522 ( .A1(n9048), .A2(n9614), .Y(n9613) );
  OR2X1_RVT U9523 ( .A1(n12295), .A2(n9615), .Y(n9609) );
  OR2X1_RVT U9524 ( .A1(n9354), .A2(n8991), .Y(n9615) );
  OR2X1_RVT U9525 ( .A1(n8974), .A2(n9000), .Y(n9608) );
  OR2X1_RVT U9526 ( .A1(n12745), .A2(n9100), .Y(n9000) );
  OR2X1_RVT U9527 ( .A1(n9474), .A2(n9388), .Y(n9597) );
  OR2X1_RVT U9528 ( .A1(n12311), .A2(n9011), .Y(n9388) );
  AND4X1_RVT U9529 ( .A1(n9617), .A2(n9618), .A3(n9619), .A4(n9620), .Y(n9616)
         );
  AND4X1_RVT U9530 ( .A1(n9621), .A2(n9622), .A3(n9623), .A4(n9624), .Y(n9620)
         );
  AND4X1_RVT U9531 ( .A1(n9625), .A2(n9626), .A3(n9627), .A4(n9628), .Y(n9624)
         );
  OR2X1_RVT U9532 ( .A1(n9462), .A2(n9606), .Y(n9628) );
  OR2X1_RVT U9533 ( .A1(n12744), .A2(n12305), .Y(n9606) );
  OR2X1_RVT U9534 ( .A1(n12279), .A2(n12289), .Y(n9462) );
  OR2X1_RVT U9535 ( .A1(n9629), .A2(n9048), .Y(n9627) );
  AND2X1_RVT U9536 ( .A1(n8994), .A2(n9561), .Y(n9629) );
  OR2X1_RVT U9537 ( .A1(n236), .A2(n9630), .Y(n8994) );
  OR2X1_RVT U9538 ( .A1(n12279), .A2(n12741), .Y(n9630) );
  OR2X1_RVT U9539 ( .A1(n9631), .A2(n8976), .Y(n9626) );
  OR2X1_RVT U9540 ( .A1(n12293), .A2(n9137), .Y(n8976) );
  AND2X1_RVT U9541 ( .A1(n9112), .A2(n9632), .Y(n9631) );
  OR2X1_RVT U9542 ( .A1(n8991), .A2(n9193), .Y(n9632) );
  OR2X1_RVT U9543 ( .A1(n12297), .A2(n12285), .Y(n8991) );
  OR2X1_RVT U9544 ( .A1(n9237), .A2(n9633), .Y(n9112) );
  OR2X1_RVT U9545 ( .A1(n12752), .A2(n12300), .Y(n9633) );
  OR2X1_RVT U9546 ( .A1(n9634), .A2(n9035), .Y(n9625) );
  AND2X1_RVT U9547 ( .A1(n9432), .A2(n9635), .Y(n9634) );
  OR2X1_RVT U9548 ( .A1(n9636), .A2(n12741), .Y(n9635) );
  AND2X1_RVT U9549 ( .A1(n9091), .A2(n9444), .Y(n9636) );
  OR2X1_RVT U9550 ( .A1(n12749), .A2(n9053), .Y(n9444) );
  OR2X1_RVT U9551 ( .A1(n12306), .A2(n9637), .Y(n9432) );
  OR2X1_RVT U9552 ( .A1(n12754), .A2(n12750), .Y(n9637) );
  OR2X1_RVT U9553 ( .A1(n9638), .A2(n12284), .Y(n9623) );
  AND2X1_RVT U9554 ( .A1(n9639), .A2(n9640), .Y(n9638) );
  OR2X1_RVT U9555 ( .A1(n9641), .A2(n9137), .Y(n9640) );
  AND2X1_RVT U9556 ( .A1(n9202), .A2(n9642), .Y(n9641) );
  OR2X1_RVT U9557 ( .A1(n8993), .A2(n9115), .Y(n9639) );
  OR2X1_RVT U9558 ( .A1(n12298), .A2(n9051), .Y(n9115) );
  OR2X1_RVT U9559 ( .A1(n9643), .A2(n12750), .Y(n9622) );
  AND2X1_RVT U9560 ( .A1(n9207), .A2(n9366), .Y(n9643) );
  OR2X1_RVT U9561 ( .A1(n12296), .A2(n9644), .Y(n9366) );
  OR2X1_RVT U9562 ( .A1(n9047), .A2(n12285), .Y(n9644) );
  OR2X1_RVT U9563 ( .A1(n8993), .A2(n9474), .Y(n9207) );
  OR2X1_RVT U9564 ( .A1(n12285), .A2(n12300), .Y(n9474) );
  OR2X1_RVT U9565 ( .A1(n9645), .A2(n12282), .Y(n9621) );
  AND2X1_RVT U9566 ( .A1(n9247), .A2(n9646), .Y(n9645) );
  OR2X1_RVT U9567 ( .A1(n9461), .A2(n9041), .Y(n9646) );
  OR2X1_RVT U9568 ( .A1(n9100), .A2(n9582), .Y(n9247) );
  OR2X1_RVT U9569 ( .A1(n12749), .A2(n236), .Y(n9582) );
  AND2X1_RVT U9570 ( .A1(n12286), .A2(n12752), .Y(n9343) );
  AND4X1_RVT U9571 ( .A1(n9647), .A2(n9648), .A3(n9649), .A4(n9650), .Y(n9619)
         );
  AND4X1_RVT U9572 ( .A1(n9651), .A2(n9652), .A3(n9653), .A4(n9654), .Y(n9650)
         );
  OR2X1_RVT U9573 ( .A1(n9655), .A2(n12291), .Y(n9654) );
  AND2X1_RVT U9574 ( .A1(n9234), .A2(n9305), .Y(n9655) );
  OR2X1_RVT U9575 ( .A1(n9050), .A2(n9561), .Y(n9305) );
  OR2X1_RVT U9576 ( .A1(n12752), .A2(n9047), .Y(n9561) );
  OR2X1_RVT U9577 ( .A1(n12739), .A2(n12281), .Y(n9050) );
  OR2X1_RVT U9578 ( .A1(n12282), .A2(n9337), .Y(n9234) );
  OR2X1_RVT U9579 ( .A1(n12286), .A2(n12300), .Y(n9337) );
  OR2X1_RVT U9580 ( .A1(n9656), .A2(n12748), .Y(n9653) );
  AND2X1_RVT U9581 ( .A1(n9396), .A2(n9657), .Y(n9656) );
  OR2X1_RVT U9582 ( .A1(n9354), .A2(n9064), .Y(n9657) );
  OR2X1_RVT U9583 ( .A1(n9237), .A2(n9658), .Y(n9064) );
  OR2X1_RVT U9584 ( .A1(n12311), .A2(n12287), .Y(n9658) );
  OR2X1_RVT U9585 ( .A1(n12295), .A2(n9659), .Y(n9396) );
  OR2X1_RVT U9586 ( .A1(n9237), .A2(n9033), .Y(n9659) );
  OR2X1_RVT U9587 ( .A1(n9660), .A2(n12754), .Y(n9652) );
  AND2X1_RVT U9588 ( .A1(n9342), .A2(n9271), .Y(n9660) );
  OR2X1_RVT U9589 ( .A1(n9053), .A2(n9089), .Y(n9271) );
  OR2X1_RVT U9590 ( .A1(n12746), .A2(n9237), .Y(n9089) );
  OR2X1_RVT U9591 ( .A1(n9461), .A2(n9069), .Y(n9342) );
  OR2X1_RVT U9592 ( .A1(n12292), .A2(n12751), .Y(n9461) );
  OR2X1_RVT U9593 ( .A1(n9661), .A2(n9111), .Y(n9651) );
  AND2X1_RVT U9594 ( .A1(n9662), .A2(n9663), .Y(n9661) );
  OR2X1_RVT U9595 ( .A1(n9033), .A2(n9460), .Y(n9663) );
  OR2X1_RVT U9596 ( .A1(n12748), .A2(n244), .Y(n9460) );
  AND2X1_RVT U9597 ( .A1(n9664), .A2(n9328), .Y(n9662) );
  OR2X1_RVT U9598 ( .A1(n9041), .A2(n9665), .Y(n9328) );
  OR2X1_RVT U9599 ( .A1(n12308), .A2(n12287), .Y(n9665) );
  OR2X1_RVT U9600 ( .A1(n9097), .A2(n9034), .Y(n9649) );
  OR2X1_RVT U9601 ( .A1(n12741), .A2(n8993), .Y(n9097) );
  OR2X1_RVT U9602 ( .A1(n9666), .A2(n8997), .Y(n9648) );
  AND2X1_RVT U9603 ( .A1(n9667), .A2(n9178), .Y(n9666) );
  AND2X1_RVT U9604 ( .A1(n9668), .A2(n9669), .Y(n9178) );
  OR2X1_RVT U9605 ( .A1(n12296), .A2(n9202), .Y(n9669) );
  OR2X1_RVT U9606 ( .A1(n9100), .A2(n8974), .Y(n9668) );
  OR2X1_RVT U9607 ( .A1(n12281), .A2(n9047), .Y(n8974) );
  AND2X1_RVT U9608 ( .A1(n9670), .A2(n9364), .Y(n9667) );
  OR2X1_RVT U9609 ( .A1(n9131), .A2(n9614), .Y(n9364) );
  OR2X1_RVT U9610 ( .A1(n12743), .A2(n234), .Y(n9614) );
  OR2X1_RVT U9611 ( .A1(n8993), .A2(n9160), .Y(n9670) );
  OR2X1_RVT U9612 ( .A1(n12280), .A2(n9671), .Y(n9160) );
  OR2X1_RVT U9613 ( .A1(n12739), .A2(n12309), .Y(n9671) );
  OR2X1_RVT U9614 ( .A1(n9672), .A2(n12739), .Y(n9647) );
  AND4X1_RVT U9615 ( .A1(n9673), .A2(n9674), .A3(n9675), .A4(n9506), .Y(n9672)
         );
  OR2X1_RVT U9616 ( .A1(n9047), .A2(n9427), .Y(n9506) );
  OR2X1_RVT U9617 ( .A1(n12744), .A2(n12750), .Y(n9427) );
  OR2X1_RVT U9618 ( .A1(n9047), .A2(n9676), .Y(n9675) );
  OR2X1_RVT U9619 ( .A1(n12286), .A2(n12291), .Y(n9676) );
  OR2X1_RVT U9620 ( .A1(n12749), .A2(n9006), .Y(n9047) );
  OR2X1_RVT U9621 ( .A1(n9677), .A2(n9128), .Y(n9674) );
  OR2X1_RVT U9622 ( .A1(n12280), .A2(n8972), .Y(n9128) );
  AND2X1_RVT U9623 ( .A1(n9111), .A2(n9678), .Y(n9677) );
  OR2X1_RVT U9624 ( .A1(n12747), .A2(n9011), .Y(n9678) );
  OR2X1_RVT U9625 ( .A1(n12743), .A2(n12291), .Y(n9111) );
  OR2X1_RVT U9626 ( .A1(n12745), .A2(n9642), .Y(n9673) );
  OR2X1_RVT U9627 ( .A1(n12749), .A2(n9051), .Y(n9642) );
  OR2X1_RVT U9628 ( .A1(n8997), .A2(n234), .Y(n9051) );
  AND4X1_RVT U9629 ( .A1(n9679), .A2(n9680), .A3(n9681), .A4(n9682), .Y(n9618)
         );
  AND4X1_RVT U9630 ( .A1(n9683), .A2(n9684), .A3(n9685), .A4(n9686), .Y(n9682)
         );
  OR2X1_RVT U9631 ( .A1(n9069), .A2(n9196), .Y(n9686) );
  OR2X1_RVT U9632 ( .A1(n12293), .A2(n9091), .Y(n9196) );
  OR2X1_RVT U9633 ( .A1(n12297), .A2(n9237), .Y(n9069) );
  OR2X1_RVT U9634 ( .A1(n9056), .A2(n9532), .Y(n9685) );
  OR2X1_RVT U9635 ( .A1(n12753), .A2(n12280), .Y(n9532) );
  OR2X1_RVT U9636 ( .A1(n9122), .A2(n9048), .Y(n9056) );
  OR2X1_RVT U9637 ( .A1(n9041), .A2(n9068), .Y(n9684) );
  OR2X1_RVT U9638 ( .A1(n12289), .A2(n12302), .Y(n9068) );
  OR2X1_RVT U9639 ( .A1(n12279), .A2(n12740), .Y(n9041) );
  OR2X1_RVT U9640 ( .A1(n244), .A2(n9407), .Y(n9683) );
  OR2X1_RVT U9641 ( .A1(n12287), .A2(n9194), .Y(n9407) );
  OR2X1_RVT U9642 ( .A1(n9011), .A2(n9441), .Y(n9681) );
  OR2X1_RVT U9643 ( .A1(n244), .A2(n9687), .Y(n9441) );
  OR2X1_RVT U9644 ( .A1(n12746), .A2(n12300), .Y(n9687) );
  AND2X1_RVT U9645 ( .A1(n12281), .A2(n12284), .Y(n9471) );
  OR2X1_RVT U9646 ( .A1(n9053), .A2(n9001), .Y(n9680) );
  OR2X1_RVT U9647 ( .A1(n12309), .A2(n9688), .Y(n9001) );
  OR2X1_RVT U9648 ( .A1(n12747), .A2(n12739), .Y(n9688) );
  OR2X1_RVT U9649 ( .A1(n12286), .A2(n9033), .Y(n9053) );
  OR2X1_RVT U9650 ( .A1(n9100), .A2(n9664), .Y(n9679) );
  OR2X1_RVT U9651 ( .A1(n12282), .A2(n9055), .Y(n9664) );
  OR2X1_RVT U9652 ( .A1(n12749), .A2(n12750), .Y(n9055) );
  AND4X1_RVT U9653 ( .A1(n9689), .A2(n9166), .A3(n9690), .A4(n9691), .Y(n9617)
         );
  OR2X1_RVT U9654 ( .A1(n12286), .A2(n9611), .Y(n9691) );
  OR2X1_RVT U9655 ( .A1(n12745), .A2(n9161), .Y(n9611) );
  OR2X1_RVT U9656 ( .A1(n12284), .A2(n9202), .Y(n9161) );
  OR2X1_RVT U9657 ( .A1(n12279), .A2(n9028), .Y(n9202) );
  AND2X1_RVT U9658 ( .A1(n9692), .A2(n9693), .Y(n9690) );
  OR2X1_RVT U9659 ( .A1(n12308), .A2(n9531), .Y(n9693) );
  OR2X1_RVT U9660 ( .A1(n9100), .A2(n9193), .Y(n9531) );
  OR2X1_RVT U9661 ( .A1(n12286), .A2(n12280), .Y(n9193) );
  OR2X1_RVT U9662 ( .A1(n12281), .A2(n8989), .Y(n9028) );
  OR2X1_RVT U9663 ( .A1(n12752), .A2(n9262), .Y(n9692) );
  OR2X1_RVT U9664 ( .A1(n12305), .A2(n9296), .Y(n9262) );
  OR2X1_RVT U9665 ( .A1(n12744), .A2(n12739), .Y(n9296) );
  OR2X1_RVT U9666 ( .A1(n12742), .A2(n12297), .Y(n8972) );
  AND2X1_RVT U9667 ( .A1(n9694), .A2(n9695), .Y(n9166) );
  OR2X1_RVT U9668 ( .A1(n9048), .A2(n9034), .Y(n9695) );
  OR2X1_RVT U9669 ( .A1(n12751), .A2(n9006), .Y(n9034) );
  AND2X1_RVT U9670 ( .A1(n9033), .A2(n8997), .Y(n9086) );
  OR2X1_RVT U9671 ( .A1(n12292), .A2(n9100), .Y(n9048) );
  OR2X1_RVT U9672 ( .A1(n12740), .A2(n9137), .Y(n9100) );
  OR2X1_RVT U9673 ( .A1(n9696), .A2(n9091), .Y(n9694) );
  OR2X1_RVT U9674 ( .A1(n12286), .A2(n234), .Y(n9091) );
  AND2X1_RVT U9675 ( .A1(n12753), .A2(n12279), .Y(n9354) );
  OR2X1_RVT U9676 ( .A1(n12285), .A2(n9194), .Y(n9696) );
  OR2X1_RVT U9677 ( .A1(n12749), .A2(n12302), .Y(n9194) );
  AND2X1_RVT U9678 ( .A1(n9697), .A2(n9698), .Y(n9689) );
  OR2X1_RVT U9679 ( .A1(n9014), .A2(n9347), .Y(n9698) );
  OR2X1_RVT U9680 ( .A1(n12287), .A2(n9054), .Y(n9347) );
  OR2X1_RVT U9681 ( .A1(n12302), .A2(n9131), .Y(n9054) );
  OR2X1_RVT U9682 ( .A1(n12282), .A2(n12285), .Y(n9131) );
  OR2X1_RVT U9683 ( .A1(n12746), .A2(n12744), .Y(n8993) );
  OR2X1_RVT U9684 ( .A1(n12754), .A2(n12748), .Y(n9014) );
  XOR2X1_RVT U9685 ( .A1(key[36]), .A2(state[36]), .Y(n8989) );
  OR2X1_RVT U9686 ( .A1(n9006), .A2(n9135), .Y(n9697) );
  OR2X1_RVT U9687 ( .A1(n9237), .A2(n9428), .Y(n9135) );
  OR2X1_RVT U9688 ( .A1(n12289), .A2(n9035), .Y(n9428) );
  OR2X1_RVT U9689 ( .A1(n12747), .A2(n9137), .Y(n9035) );
  XOR2X1_RVT U9690 ( .A1(key[34]), .A2(state[34]), .Y(n9137) );
  XOR2X1_RVT U9691 ( .A1(key[35]), .A2(state[35]), .Y(n9071) );
  OR2X1_RVT U9692 ( .A1(n12752), .A2(n12287), .Y(n9011) );
  XOR2X1_RVT U9693 ( .A1(key[37]), .A2(state[37]), .Y(n8997) );
  XOR2X1_RVT U9694 ( .A1(key[38]), .A2(state[38]), .Y(n9033) );
  OR2X1_RVT U9695 ( .A1(n12742), .A2(n12285), .Y(n9237) );
  XOR2X1_RVT U9696 ( .A1(key[32]), .A2(state[32]), .Y(n9012) );
  XOR2X1_RVT U9697 ( .A1(key[33]), .A2(state[33]), .Y(n9122) );
  XOR2X1_RVT U9698 ( .A1(key[39]), .A2(state[39]), .Y(n9006) );
  AND4X1_RVT U9699 ( .A1(n9700), .A2(n9701), .A3(n9702), .A4(n9703), .Y(n9699)
         );
  AND4X1_RVT U9700 ( .A1(n9704), .A2(n9705), .A3(n9706), .A4(n9707), .Y(n9703)
         );
  AND4X1_RVT U9701 ( .A1(n9708), .A2(n9709), .A3(n9710), .A4(n9711), .Y(n9707)
         );
  OR2X1_RVT U9702 ( .A1(n12273), .A2(n9713), .Y(n9706) );
  OR2X1_RVT U9703 ( .A1(n9714), .A2(n9715), .Y(n9704) );
  OR2X1_RVT U9704 ( .A1(n12864), .A2(n9716), .Y(n9715) );
  AND4X1_RVT U9705 ( .A1(n9717), .A2(n9718), .A3(n9719), .A4(n9720), .Y(n9702)
         );
  OR2X1_RVT U9706 ( .A1(n9721), .A2(n12862), .Y(n9720) );
  AND2X1_RVT U9707 ( .A1(n9722), .A2(n9723), .Y(n9721) );
  AND2X1_RVT U9708 ( .A1(n9724), .A2(n9725), .Y(n9719) );
  OR2X1_RVT U9709 ( .A1(n9726), .A2(n96), .Y(n9725) );
  AND2X1_RVT U9710 ( .A1(n9727), .A2(n9728), .Y(n9726) );
  OR2X1_RVT U9711 ( .A1(n12264), .A2(n9730), .Y(n9728) );
  OR2X1_RVT U9712 ( .A1(n9716), .A2(n9731), .Y(n9727) );
  OR2X1_RVT U9713 ( .A1(n9732), .A2(n12270), .Y(n9724) );
  AND2X1_RVT U9714 ( .A1(n9734), .A2(n9735), .Y(n9732) );
  OR2X1_RVT U9715 ( .A1(n9736), .A2(n9737), .Y(n9718) );
  AND2X1_RVT U9716 ( .A1(n9738), .A2(n9739), .Y(n9736) );
  OR2X1_RVT U9717 ( .A1(n12265), .A2(n9740), .Y(n9739) );
  AND2X1_RVT U9718 ( .A1(n9741), .A2(n9742), .Y(n9738) );
  AND2X1_RVT U9719 ( .A1(n9743), .A2(n9744), .Y(n9717) );
  OR2X1_RVT U9720 ( .A1(n9745), .A2(n12247), .Y(n9744) );
  AND2X1_RVT U9721 ( .A1(n9747), .A2(n9748), .Y(n9745) );
  OR2X1_RVT U9722 ( .A1(n9749), .A2(n9750), .Y(n9748) );
  OR2X1_RVT U9723 ( .A1(n12256), .A2(n12251), .Y(n9750) );
  OR2X1_RVT U9724 ( .A1(n9753), .A2(n9754), .Y(n9743) );
  AND2X1_RVT U9725 ( .A1(n9755), .A2(n9756), .Y(n9753) );
  AND2X1_RVT U9726 ( .A1(n9757), .A2(n9758), .Y(n9755) );
  AND4X1_RVT U9727 ( .A1(n9759), .A2(n9760), .A3(n9761), .A4(n9762), .Y(n9701)
         );
  AND4X1_RVT U9728 ( .A1(n9763), .A2(n9764), .A3(n9765), .A4(n9766), .Y(n9762)
         );
  OR2X1_RVT U9729 ( .A1(n9767), .A2(n12276), .Y(n9766) );
  AND4X1_RVT U9730 ( .A1(n9769), .A2(n9770), .A3(n9771), .A4(n9772), .Y(n9767)
         );
  OR2X1_RVT U9731 ( .A1(n9773), .A2(n9740), .Y(n9772) );
  OR2X1_RVT U9732 ( .A1(n9774), .A2(n12262), .Y(n9771) );
  OR2X1_RVT U9733 ( .A1(n9776), .A2(n12253), .Y(n9765) );
  AND4X1_RVT U9734 ( .A1(n9777), .A2(n9778), .A3(n9779), .A4(n9780), .Y(n9776)
         );
  OR2X1_RVT U9735 ( .A1(n9781), .A2(n9782), .Y(n9780) );
  OR2X1_RVT U9736 ( .A1(n12270), .A2(n12265), .Y(n9782) );
  AND2X1_RVT U9737 ( .A1(n9783), .A2(n9784), .Y(n9779) );
  OR2X1_RVT U9738 ( .A1(n12866), .A2(n9785), .Y(n9778) );
  OR2X1_RVT U9739 ( .A1(n9786), .A2(n9787), .Y(n9777) );
  AND2X1_RVT U9740 ( .A1(n9788), .A2(n9789), .Y(n9786) );
  OR2X1_RVT U9741 ( .A1(n12270), .A2(n9790), .Y(n9789) );
  OR2X1_RVT U9742 ( .A1(n9723), .A2(n9791), .Y(n9764) );
  OR2X1_RVT U9743 ( .A1(n9790), .A2(n9792), .Y(n9763) );
  OR2X1_RVT U9744 ( .A1(n9793), .A2(n9794), .Y(n9761) );
  OR2X1_RVT U9745 ( .A1(n9795), .A2(n9788), .Y(n9760) );
  OR2X1_RVT U9746 ( .A1(n9796), .A2(n9797), .Y(n9759) );
  AND4X1_RVT U9747 ( .A1(n9798), .A2(n9799), .A3(n9800), .A4(n9801), .Y(n9700)
         );
  AND2X1_RVT U9748 ( .A1(n9802), .A2(n9803), .Y(n9801) );
  OR2X1_RVT U9749 ( .A1(n9787), .A2(n9804), .Y(n9803) );
  AND2X1_RVT U9750 ( .A1(n9805), .A2(n9806), .Y(n9802) );
  OR2X1_RVT U9751 ( .A1(n9807), .A2(n9730), .Y(n9806) );
  OR2X1_RVT U9752 ( .A1(n9731), .A2(n9808), .Y(n9805) );
  OR2X1_RVT U9753 ( .A1(n94), .A2(n9809), .Y(n9800) );
  OR2X1_RVT U9754 ( .A1(n9810), .A2(n12260), .Y(n9799) );
  OR2X1_RVT U9755 ( .A1(n12263), .A2(n9812), .Y(n9798) );
  AND4X1_RVT U9756 ( .A1(n9814), .A2(n9815), .A3(n9816), .A4(n9817), .Y(n9813)
         );
  AND4X1_RVT U9757 ( .A1(n9818), .A2(n9709), .A3(n9819), .A4(n9820), .Y(n9817)
         );
  AND4X1_RVT U9758 ( .A1(n9821), .A2(n9822), .A3(n9823), .A4(n9824), .Y(n9820)
         );
  OR2X1_RVT U9759 ( .A1(n9730), .A2(n9825), .Y(n9824) );
  OR2X1_RVT U9760 ( .A1(n9826), .A2(n12275), .Y(n9825) );
  OR2X1_RVT U9761 ( .A1(n9731), .A2(n9827), .Y(n9823) );
  OR2X1_RVT U9762 ( .A1(n94), .A2(n12259), .Y(n9827) );
  OR2X1_RVT U9763 ( .A1(n9828), .A2(n9774), .Y(n9822) );
  AND2X1_RVT U9764 ( .A1(n9785), .A2(n9829), .Y(n9828) );
  OR2X1_RVT U9765 ( .A1(n9830), .A2(n9831), .Y(n9821) );
  AND2X1_RVT U9766 ( .A1(n9832), .A2(n9833), .Y(n9830) );
  AND2X1_RVT U9767 ( .A1(n9834), .A2(n9835), .Y(n9819) );
  OR2X1_RVT U9768 ( .A1(n9781), .A2(n9836), .Y(n9835) );
  OR2X1_RVT U9769 ( .A1(n9837), .A2(n12864), .Y(n9836) );
  OR2X1_RVT U9770 ( .A1(n9838), .A2(n9839), .Y(n9834) );
  OR2X1_RVT U9771 ( .A1(n9840), .A2(n12264), .Y(n9839) );
  OR2X1_RVT U9772 ( .A1(n9716), .A2(n9841), .Y(n9709) );
  AND4X1_RVT U9773 ( .A1(n9842), .A2(n9843), .A3(n9844), .A4(n9845), .Y(n9816)
         );
  AND4X1_RVT U9774 ( .A1(n9846), .A2(n9847), .A3(n9848), .A4(n9849), .Y(n9845)
         );
  OR2X1_RVT U9775 ( .A1(n9850), .A2(n12278), .Y(n9849) );
  AND2X1_RVT U9776 ( .A1(n9852), .A2(n9853), .Y(n9850) );
  OR2X1_RVT U9777 ( .A1(n12247), .A2(n9731), .Y(n9853) );
  OR2X1_RVT U9778 ( .A1(n9854), .A2(n9733), .Y(n9848) );
  AND2X1_RVT U9779 ( .A1(n9855), .A2(n9856), .Y(n9854) );
  OR2X1_RVT U9780 ( .A1(n9857), .A2(n12863), .Y(n9847) );
  AND2X1_RVT U9781 ( .A1(n9858), .A2(n9859), .Y(n9857) );
  OR2X1_RVT U9782 ( .A1(n9860), .A2(n9809), .Y(n9859) );
  AND2X1_RVT U9783 ( .A1(n12278), .A2(n12262), .Y(n9860) );
  OR2X1_RVT U9784 ( .A1(n9861), .A2(n12248), .Y(n9846) );
  AND2X1_RVT U9785 ( .A1(n9863), .A2(n9864), .Y(n9861) );
  OR2X1_RVT U9786 ( .A1(n9865), .A2(n12254), .Y(n9844) );
  AND2X1_RVT U9787 ( .A1(n9866), .A2(n9867), .Y(n9865) );
  OR2X1_RVT U9788 ( .A1(n12262), .A2(n9868), .Y(n9867) );
  AND2X1_RVT U9789 ( .A1(n9869), .A2(n9870), .Y(n9866) );
  OR2X1_RVT U9790 ( .A1(n9871), .A2(n9872), .Y(n9869) );
  OR2X1_RVT U9791 ( .A1(n9716), .A2(n9787), .Y(n9872) );
  OR2X1_RVT U9792 ( .A1(n9873), .A2(n12860), .Y(n9843) );
  AND2X1_RVT U9793 ( .A1(n9874), .A2(n9875), .Y(n9873) );
  OR2X1_RVT U9794 ( .A1(n9876), .A2(n9877), .Y(n9842) );
  AND2X1_RVT U9795 ( .A1(n9878), .A2(n9879), .Y(n9876) );
  AND2X1_RVT U9796 ( .A1(n9880), .A2(n9881), .Y(n9878) );
  OR2X1_RVT U9797 ( .A1(n96), .A2(n9809), .Y(n9881) );
  OR2X1_RVT U9798 ( .A1(n12272), .A2(n9774), .Y(n9880) );
  AND4X1_RVT U9799 ( .A1(n9882), .A2(n9883), .A3(n9884), .A4(n9885), .Y(n9815)
         );
  AND4X1_RVT U9800 ( .A1(n9886), .A2(n9887), .A3(n9888), .A4(n9889), .Y(n9885)
         );
  OR2X1_RVT U9801 ( .A1(n9809), .A2(n9808), .Y(n9889) );
  OR2X1_RVT U9802 ( .A1(n9740), .A2(n9890), .Y(n9888) );
  OR2X1_RVT U9803 ( .A1(n9773), .A2(n9891), .Y(n9887) );
  OR2X1_RVT U9804 ( .A1(n9716), .A2(n9892), .Y(n9886) );
  AND2X1_RVT U9805 ( .A1(n9893), .A2(n9894), .Y(n9884) );
  OR2X1_RVT U9806 ( .A1(n12273), .A2(n9895), .Y(n9894) );
  OR2X1_RVT U9807 ( .A1(n12252), .A2(n9792), .Y(n9893) );
  OR2X1_RVT U9808 ( .A1(n9896), .A2(n9751), .Y(n9883) );
  AND4X1_RVT U9809 ( .A1(n9897), .A2(n9898), .A3(n9899), .A4(n9900), .Y(n9896)
         );
  OR2X1_RVT U9810 ( .A1(n9901), .A2(n9716), .Y(n9899) );
  OR2X1_RVT U9811 ( .A1(n12852), .A2(n9902), .Y(n9898) );
  OR2X1_RVT U9812 ( .A1(n9903), .A2(n12860), .Y(n9897) );
  AND2X1_RVT U9813 ( .A1(n9794), .A2(n9904), .Y(n9903) );
  OR2X1_RVT U9814 ( .A1(n9796), .A2(n9905), .Y(n9882) );
  AND4X1_RVT U9815 ( .A1(n9906), .A2(n9907), .A3(n9908), .A4(n9909), .Y(n9814)
         );
  AND4X1_RVT U9816 ( .A1(n9910), .A2(n9911), .A3(n9912), .A4(n9913), .Y(n9909)
         );
  OR2X1_RVT U9817 ( .A1(n12856), .A2(n9914), .Y(n9913) );
  OR2X1_RVT U9818 ( .A1(n12857), .A2(n9915), .Y(n9912) );
  OR2X1_RVT U9819 ( .A1(n12854), .A2(n9916), .Y(n9911) );
  OR2X1_RVT U9820 ( .A1(n12246), .A2(n9917), .Y(n9910) );
  OR2X1_RVT U9821 ( .A1(n9918), .A2(n12253), .Y(n9907) );
  AND4X1_RVT U9822 ( .A1(n9920), .A2(n9921), .A3(n9922), .A4(n9923), .Y(n9919)
         );
  AND4X1_RVT U9823 ( .A1(n9924), .A2(n9925), .A3(n9926), .A4(n9927), .Y(n9923)
         );
  AND4X1_RVT U9824 ( .A1(n9928), .A2(n9705), .A3(n9875), .A4(n9929), .Y(n9927)
         );
  OR2X1_RVT U9825 ( .A1(n9930), .A2(n12851), .Y(n9705) );
  AND2X1_RVT U9826 ( .A1(n9931), .A2(n9932), .Y(n9930) );
  OR2X1_RVT U9827 ( .A1(n9749), .A2(n9933), .Y(n9932) );
  OR2X1_RVT U9828 ( .A1(n9934), .A2(n9831), .Y(n9931) );
  OR2X1_RVT U9829 ( .A1(n9935), .A2(n9790), .Y(n9928) );
  AND2X1_RVT U9830 ( .A1(n9936), .A2(n9937), .Y(n9935) );
  OR2X1_RVT U9831 ( .A1(n12856), .A2(n9774), .Y(n9937) );
  OR2X1_RVT U9832 ( .A1(n9938), .A2(n9733), .Y(n9926) );
  AND2X1_RVT U9833 ( .A1(n9939), .A2(n9940), .Y(n9938) );
  OR2X1_RVT U9834 ( .A1(n9941), .A2(n12862), .Y(n9940) );
  AND2X1_RVT U9835 ( .A1(n9781), .A2(n9942), .Y(n9941) );
  OR2X1_RVT U9836 ( .A1(n9943), .A2(n12273), .Y(n9925) );
  AND2X1_RVT U9837 ( .A1(n9944), .A2(n9945), .Y(n9943) );
  OR2X1_RVT U9838 ( .A1(n9774), .A2(n9740), .Y(n9945) );
  OR2X1_RVT U9839 ( .A1(n9946), .A2(n12256), .Y(n9924) );
  AND2X1_RVT U9840 ( .A1(n9858), .A2(n9947), .Y(n9946) );
  OR2X1_RVT U9841 ( .A1(n9787), .A2(n9948), .Y(n9858) );
  AND4X1_RVT U9842 ( .A1(n9949), .A2(n9950), .A3(n9951), .A4(n9952), .Y(n9922)
         );
  OR2X1_RVT U9843 ( .A1(n9953), .A2(n12263), .Y(n9952) );
  AND2X1_RVT U9844 ( .A1(n9954), .A2(n9955), .Y(n9953) );
  OR2X1_RVT U9845 ( .A1(n9831), .A2(n9731), .Y(n9955) );
  AND2X1_RVT U9846 ( .A1(n9956), .A2(n9957), .Y(n9954) );
  OR2X1_RVT U9847 ( .A1(n9871), .A2(n9933), .Y(n9956) );
  AND2X1_RVT U9848 ( .A1(n9958), .A2(n9959), .Y(n9951) );
  OR2X1_RVT U9849 ( .A1(n9960), .A2(n9862), .Y(n9959) );
  AND2X1_RVT U9850 ( .A1(n9961), .A2(n9770), .Y(n9960) );
  OR2X1_RVT U9851 ( .A1(n9716), .A2(n9831), .Y(n9770) );
  OR2X1_RVT U9852 ( .A1(n9962), .A2(n96), .Y(n9958) );
  AND2X1_RVT U9853 ( .A1(n9963), .A2(n9964), .Y(n9962) );
  OR2X1_RVT U9854 ( .A1(n9965), .A2(n12265), .Y(n9964) );
  AND2X1_RVT U9855 ( .A1(n9966), .A2(n9967), .Y(n9965) );
  OR2X1_RVT U9856 ( .A1(n12260), .A2(n9781), .Y(n9967) );
  OR2X1_RVT U9857 ( .A1(n12866), .A2(n12262), .Y(n9966) );
  AND2X1_RVT U9858 ( .A1(n9832), .A2(n9942), .Y(n9963) );
  OR2X1_RVT U9859 ( .A1(n9862), .A2(n9968), .Y(n9832) );
  OR2X1_RVT U9860 ( .A1(n12861), .A2(n12857), .Y(n9968) );
  OR2X1_RVT U9861 ( .A1(n9969), .A2(n9851), .Y(n9950) );
  AND4X1_RVT U9862 ( .A1(n9810), .A2(n9970), .A3(n9971), .A4(n9972), .Y(n9969)
         );
  OR2X1_RVT U9863 ( .A1(n12264), .A2(n9831), .Y(n9972) );
  AND2X1_RVT U9864 ( .A1(n9973), .A2(n9974), .Y(n9971) );
  OR2X1_RVT U9865 ( .A1(n12866), .A2(n12273), .Y(n9970) );
  AND2X1_RVT U9866 ( .A1(n9975), .A2(n9976), .Y(n9810) );
  OR2X1_RVT U9867 ( .A1(n9977), .A2(n94), .Y(n9976) );
  OR2X1_RVT U9868 ( .A1(n9774), .A2(n12851), .Y(n9975) );
  AND2X1_RVT U9869 ( .A1(n9978), .A2(n9979), .Y(n9949) );
  OR2X1_RVT U9870 ( .A1(n9980), .A2(n12853), .Y(n9979) );
  AND2X1_RVT U9871 ( .A1(n9981), .A2(n9982), .Y(n9980) );
  OR2X1_RVT U9872 ( .A1(n9983), .A2(n12267), .Y(n9982) );
  AND2X1_RVT U9873 ( .A1(n9984), .A2(n9985), .Y(n9983) );
  AND2X1_RVT U9874 ( .A1(n9986), .A2(n9987), .Y(n9981) );
  OR2X1_RVT U9875 ( .A1(n9988), .A2(n12276), .Y(n9978) );
  AND4X1_RVT U9876 ( .A1(n9989), .A2(n9990), .A3(n9991), .A4(n9992), .Y(n9988)
         );
  OR2X1_RVT U9877 ( .A1(n12865), .A2(n9993), .Y(n9991) );
  OR2X1_RVT U9878 ( .A1(n94), .A2(n9788), .Y(n9990) );
  OR2X1_RVT U9879 ( .A1(n9877), .A2(n9831), .Y(n9989) );
  AND4X1_RVT U9880 ( .A1(n9994), .A2(n9995), .A3(n9996), .A4(n9997), .Y(n9921)
         );
  AND2X1_RVT U9881 ( .A1(n9998), .A2(n9841), .Y(n9997) );
  OR2X1_RVT U9882 ( .A1(n12251), .A2(n9807), .Y(n9841) );
  AND2X1_RVT U9883 ( .A1(n9999), .A2(n10000), .Y(n9998) );
  OR2X1_RVT U9884 ( .A1(n10001), .A2(n9756), .Y(n10000) );
  OR2X1_RVT U9885 ( .A1(n9808), .A2(n9868), .Y(n9999) );
  OR2X1_RVT U9886 ( .A1(n94), .A2(n10002), .Y(n9996) );
  OR2X1_RVT U9887 ( .A1(n12864), .A2(n10003), .Y(n9995) );
  OR2X1_RVT U9888 ( .A1(n9877), .A2(n10004), .Y(n9994) );
  AND4X1_RVT U9889 ( .A1(n10005), .A2(n10006), .A3(n10007), .A4(n10008), .Y(
        n9920) );
  AND2X1_RVT U9890 ( .A1(n10009), .A2(n10010), .Y(n10008) );
  OR2X1_RVT U9891 ( .A1(n12246), .A2(n10011), .Y(n10010) );
  AND2X1_RVT U9892 ( .A1(n10012), .A2(n10013), .Y(n10009) );
  OR2X1_RVT U9893 ( .A1(n9773), .A2(n9783), .Y(n10013) );
  OR2X1_RVT U9894 ( .A1(n12267), .A2(n9833), .Y(n9783) );
  OR2X1_RVT U9895 ( .A1(n12253), .A2(n10014), .Y(n10012) );
  OR2X1_RVT U9896 ( .A1(n9754), .A2(n9747), .Y(n10007) );
  OR2X1_RVT U9897 ( .A1(n9840), .A2(n10015), .Y(n9747) );
  OR2X1_RVT U9898 ( .A1(n12860), .A2(n10016), .Y(n10006) );
  OR2X1_RVT U9899 ( .A1(n12265), .A2(n9874), .Y(n10005) );
  OR2X1_RVT U9900 ( .A1(n12851), .A2(n9936), .Y(n9874) );
  AND4X1_RVT U9901 ( .A1(n10018), .A2(n10019), .A3(n10020), .A4(n10021), .Y(
        n10017) );
  AND4X1_RVT U9902 ( .A1(n10022), .A2(n10023), .A3(n10024), .A4(n10025), .Y(
        n10021) );
  AND4X1_RVT U9903 ( .A1(n10026), .A2(n10027), .A3(n6125), .A4(n10028), .Y(
        n10025) );
  OR2X1_RVT U9904 ( .A1(n8127), .A2(n10029), .Y(n6125) );
  OR2X1_RVT U9905 ( .A1(n12208), .A2(n12203), .Y(n10029) );
  OR2X1_RVT U9906 ( .A1(n12868), .A2(n72), .Y(n8127) );
  OR2X1_RVT U9907 ( .A1(n10030), .A2(n12926), .Y(n10027) );
  AND2X1_RVT U9908 ( .A1(n6208), .A2(n10031), .Y(n10030) );
  OR2X1_RVT U9909 ( .A1(n10032), .A2(n12875), .Y(n10031) );
  AND2X1_RVT U9910 ( .A1(n12201), .A2(n83), .Y(n10032) );
  OR2X1_RVT U9911 ( .A1(n12867), .A2(n8121), .Y(n6208) );
  OR2X1_RVT U9912 ( .A1(n10033), .A2(n12203), .Y(n10026) );
  AND2X1_RVT U9913 ( .A1(n1400), .A2(n10034), .Y(n10033) );
  OR2X1_RVT U9914 ( .A1(n8919), .A2(n1391), .Y(n10034) );
  OR2X1_RVT U9915 ( .A1(n12876), .A2(n7007), .Y(n1400) );
  OR2X1_RVT U9916 ( .A1(n12191), .A2(n76), .Y(n7007) );
  OR2X1_RVT U9917 ( .A1(n10035), .A2(n76), .Y(n10024) );
  AND2X1_RVT U9918 ( .A1(n10036), .A2(n10037), .Y(n10035) );
  OR2X1_RVT U9919 ( .A1(n7034), .A2(n1329), .Y(n10037) );
  AND2X1_RVT U9920 ( .A1(n8121), .A2(n8077), .Y(n10036) );
  OR2X1_RVT U9921 ( .A1(n12199), .A2(n10038), .Y(n8077) );
  OR2X1_RVT U9922 ( .A1(n71), .A2(n1312), .Y(n10038) );
  OR2X1_RVT U9923 ( .A1(n12212), .A2(n72), .Y(n8121) );
  OR2X1_RVT U9924 ( .A1(n10039), .A2(n12871), .Y(n10023) );
  AND2X1_RVT U9925 ( .A1(n7015), .A2(n8955), .Y(n10039) );
  OR2X1_RVT U9926 ( .A1(n12208), .A2(n1329), .Y(n8955) );
  OR2X1_RVT U9927 ( .A1(n69), .A2(n1370), .Y(n7015) );
  OR2X1_RVT U9928 ( .A1(n10040), .A2(n1350), .Y(n10022) );
  AND2X1_RVT U9929 ( .A1(n1389), .A2(n10041), .Y(n10040) );
  OR2X1_RVT U9930 ( .A1(n6198), .A2(n7030), .Y(n10041) );
  OR2X1_RVT U9931 ( .A1(n12212), .A2(n10042), .Y(n1389) );
  AND4X1_RVT U9932 ( .A1(n10043), .A2(n10044), .A3(n10045), .A4(n10046), .Y(
        n10020) );
  AND4X1_RVT U9933 ( .A1(n10047), .A2(n10048), .A3(n10049), .A4(n10050), .Y(
        n10046) );
  OR2X1_RVT U9934 ( .A1(n10051), .A2(n12201), .Y(n10050) );
  AND2X1_RVT U9935 ( .A1(n10052), .A2(n10053), .Y(n10051) );
  OR2X1_RVT U9936 ( .A1(n12208), .A2(n10054), .Y(n10053) );
  OR2X1_RVT U9937 ( .A1(n12874), .A2(n12867), .Y(n10054) );
  AND2X1_RVT U9938 ( .A1(n6205), .A2(n10055), .Y(n10052) );
  OR2X1_RVT U9939 ( .A1(n73), .A2(n10056), .Y(n6205) );
  OR2X1_RVT U9940 ( .A1(n10057), .A2(n1356), .Y(n10049) );
  AND2X1_RVT U9941 ( .A1(n10058), .A2(n7013), .Y(n10057) );
  AND2X1_RVT U9942 ( .A1(n6213), .A2(n1321), .Y(n10058) );
  OR2X1_RVT U9943 ( .A1(n1391), .A2(n10059), .Y(n1321) );
  OR2X1_RVT U9944 ( .A1(n12149), .A2(n1312), .Y(n10059) );
  OR2X1_RVT U9945 ( .A1(n12877), .A2(n7052), .Y(n6213) );
  OR2X1_RVT U9946 ( .A1(n10060), .A2(n12186), .Y(n10048) );
  AND2X1_RVT U9947 ( .A1(n10061), .A2(n10062), .Y(n10060) );
  OR2X1_RVT U9948 ( .A1(n10063), .A2(n12196), .Y(n10047) );
  AND4X1_RVT U9949 ( .A1(n10064), .A2(n10065), .A3(n6963), .A4(n7042), .Y(
        n10063) );
  OR2X1_RVT U9950 ( .A1(n12192), .A2(n1346), .Y(n7042) );
  OR2X1_RVT U9951 ( .A1(n1391), .A2(n8946), .Y(n6963) );
  OR2X1_RVT U9952 ( .A1(n8063), .A2(n1348), .Y(n10065) );
  OR2X1_RVT U9953 ( .A1(n10066), .A2(n12199), .Y(n10064) );
  AND2X1_RVT U9954 ( .A1(n10067), .A2(n10068), .Y(n10066) );
  OR2X1_RVT U9955 ( .A1(n71), .A2(n12875), .Y(n10068) );
  OR2X1_RVT U9956 ( .A1(n12871), .A2(n1312), .Y(n10067) );
  OR2X1_RVT U9957 ( .A1(n6190), .A2(n10056), .Y(n10045) );
  OR2X1_RVT U9958 ( .A1(n10069), .A2(n12189), .Y(n10044) );
  AND4X1_RVT U9959 ( .A1(n10070), .A2(n10071), .A3(n10072), .A4(n6964), .Y(
        n10069) );
  OR2X1_RVT U9960 ( .A1(n1323), .A2(n10073), .Y(n6964) );
  AND2X1_RVT U9961 ( .A1(n6175), .A2(n1358), .Y(n10072) );
  OR2X1_RVT U9962 ( .A1(n69), .A2(n6143), .Y(n1358) );
  OR2X1_RVT U9963 ( .A1(n12206), .A2(n10074), .Y(n6175) );
  OR2X1_RVT U9964 ( .A1(n83), .A2(n12195), .Y(n10074) );
  OR2X1_RVT U9965 ( .A1(n1314), .A2(n10075), .Y(n10070) );
  OR2X1_RVT U9966 ( .A1(n8919), .A2(n12199), .Y(n10075) );
  OR2X1_RVT U9967 ( .A1(n1325), .A2(n8917), .Y(n10043) );
  AND4X1_RVT U9968 ( .A1(n10076), .A2(n10077), .A3(n10078), .A4(n10079), .Y(
        n10019) );
  AND4X1_RVT U9969 ( .A1(n10080), .A2(n10081), .A3(n10082), .A4(n10083), .Y(
        n10079) );
  OR2X1_RVT U9970 ( .A1(n8088), .A2(n6198), .Y(n10083) );
  OR2X1_RVT U9971 ( .A1(n10073), .A2(n7000), .Y(n10082) );
  OR2X1_RVT U9972 ( .A1(n12872), .A2(n12206), .Y(n7000) );
  OR2X1_RVT U9973 ( .A1(n1323), .A2(n10084), .Y(n10081) );
  OR2X1_RVT U9974 ( .A1(n1359), .A2(n1388), .Y(n10080) );
  OR2X1_RVT U9975 ( .A1(n12188), .A2(n6198), .Y(n1359) );
  OR2X1_RVT U9976 ( .A1(n73), .A2(n7031), .Y(n10078) );
  OR2X1_RVT U9977 ( .A1(n6145), .A2(n1348), .Y(n10077) );
  OR2X1_RVT U9978 ( .A1(n8055), .A2(n12189), .Y(n1348) );
  OR2X1_RVT U9979 ( .A1(n71), .A2(n8053), .Y(n10076) );
  OR2X1_RVT U9980 ( .A1(n78), .A2(n10085), .Y(n8053) );
  OR2X1_RVT U9981 ( .A1(n12869), .A2(n72), .Y(n10085) );
  AND4X1_RVT U9982 ( .A1(n10086), .A2(n10087), .A3(n10088), .A4(n10089), .Y(
        n10018) );
  AND4X1_RVT U9983 ( .A1(n10090), .A2(n10091), .A3(n10092), .A4(n10093), .Y(
        n10089) );
  OR2X1_RVT U9984 ( .A1(n12149), .A2(n8954), .Y(n10093) );
  OR2X1_RVT U9985 ( .A1(n12871), .A2(n1306), .Y(n8954) );
  OR2X1_RVT U9986 ( .A1(n12868), .A2(n1317), .Y(n10092) );
  OR2X1_RVT U9987 ( .A1(n6145), .A2(n1386), .Y(n1317) );
  OR2X1_RVT U9988 ( .A1(n12191), .A2(n8935), .Y(n10091) );
  OR2X1_RVT U9989 ( .A1(n12186), .A2(n6989), .Y(n8935) );
  OR2X1_RVT U9990 ( .A1(n8063), .A2(n10094), .Y(n10090) );
  OR2X1_RVT U9991 ( .A1(n12873), .A2(n10095), .Y(n10088) );
  OR2X1_RVT U9992 ( .A1(n6197), .A2(n8890), .Y(n10087) );
  OR2X1_RVT U9993 ( .A1(n12190), .A2(n12184), .Y(n8890) );
  OR2X1_RVT U9994 ( .A1(n83), .A2(n1319), .Y(n10086) );
  OR2X1_RVT U9995 ( .A1(n79), .A2(n1365), .Y(n1319) );
  AND2X1_RVT U9996 ( .A1(n12188), .A2(n12196), .Y(n6131) );
  AND4X1_RVT U9997 ( .A1(n10097), .A2(n10098), .A3(n10099), .A4(n10100), .Y(
        n10096) );
  AND4X1_RVT U9998 ( .A1(n10101), .A2(n10102), .A3(n10103), .A4(n10104), .Y(
        n10100) );
  OR2X1_RVT U9999 ( .A1(n104), .A2(n10105), .Y(n10104) );
  OR2X1_RVT U10000 ( .A1(n10106), .A2(n12278), .Y(n10105) );
  AND2X1_RVT U10001 ( .A1(n12267), .A2(n9793), .Y(n10106) );
  AND2X1_RVT U10002 ( .A1(n9708), .A2(n10107), .Y(n10103) );
  OR2X1_RVT U10003 ( .A1(n12256), .A2(n10108), .Y(n9708) );
  OR2X1_RVT U10004 ( .A1(n104), .A2(n9787), .Y(n10108) );
  OR2X1_RVT U10005 ( .A1(n10109), .A2(n9716), .Y(n10102) );
  AND2X1_RVT U10006 ( .A1(n10110), .A2(n10111), .Y(n10109) );
  AND2X1_RVT U10007 ( .A1(n10112), .A2(n10113), .Y(n10101) );
  OR2X1_RVT U10008 ( .A1(n10114), .A2(n10115), .Y(n10113) );
  AND2X1_RVT U10009 ( .A1(n10116), .A2(n9797), .Y(n10114) );
  OR2X1_RVT U10010 ( .A1(n10117), .A2(n9788), .Y(n10112) );
  AND2X1_RVT U10011 ( .A1(n9973), .A2(n9807), .Y(n10117) );
  OR2X1_RVT U10012 ( .A1(n12254), .A2(n10118), .Y(n9973) );
  OR2X1_RVT U10013 ( .A1(n12866), .A2(n12264), .Y(n10118) );
  AND4X1_RVT U10014 ( .A1(n10119), .A2(n10120), .A3(n10121), .A4(n10122), .Y(
        n10099) );
  OR2X1_RVT U10015 ( .A1(n10123), .A2(n12856), .Y(n10122) );
  AND2X1_RVT U10016 ( .A1(n9856), .A2(n10124), .Y(n10123) );
  OR2X1_RVT U10017 ( .A1(n12864), .A2(n9901), .Y(n9856) );
  AND2X1_RVT U10018 ( .A1(n10125), .A2(n10126), .Y(n10121) );
  OR2X1_RVT U10019 ( .A1(n10127), .A2(n12854), .Y(n10126) );
  AND2X1_RVT U10020 ( .A1(n10128), .A2(n10129), .Y(n10127) );
  OR2X1_RVT U10021 ( .A1(n9751), .A2(n9993), .Y(n10129) );
  OR2X1_RVT U10022 ( .A1(n10130), .A2(n12852), .Y(n10125) );
  AND2X1_RVT U10023 ( .A1(n10131), .A2(n10132), .Y(n10130) );
  OR2X1_RVT U10024 ( .A1(n10133), .A2(n12267), .Y(n10120) );
  AND2X1_RVT U10025 ( .A1(n10134), .A2(n10135), .Y(n10133) );
  AND2X1_RVT U10026 ( .A1(n10136), .A2(n10137), .Y(n10134) );
  AND2X1_RVT U10027 ( .A1(n10138), .A2(n10139), .Y(n10119) );
  OR2X1_RVT U10028 ( .A1(n10140), .A2(n9977), .Y(n10139) );
  AND2X1_RVT U10029 ( .A1(n10141), .A2(n9808), .Y(n10140) );
  AND2X1_RVT U10030 ( .A1(n10142), .A2(n10143), .Y(n10141) );
  OR2X1_RVT U10031 ( .A1(n10144), .A2(n12270), .Y(n10138) );
  AND2X1_RVT U10032 ( .A1(n10145), .A2(n10146), .Y(n10144) );
  OR2X1_RVT U10033 ( .A1(n12863), .A2(n12272), .Y(n10146) );
  AND2X1_RVT U10034 ( .A1(n9797), .A2(n10147), .Y(n10145) );
  AND4X1_RVT U10035 ( .A1(n10148), .A2(n10149), .A3(n10150), .A4(n10151), .Y(
        n10098) );
  AND2X1_RVT U10036 ( .A1(n10152), .A2(n10153), .Y(n10151) );
  OR2X1_RVT U10037 ( .A1(n9790), .A2(n9864), .Y(n10153) );
  OR2X1_RVT U10038 ( .A1(n12858), .A2(n9797), .Y(n9864) );
  AND2X1_RVT U10039 ( .A1(n10154), .A2(n10155), .Y(n10152) );
  OR2X1_RVT U10040 ( .A1(n9942), .A2(n9756), .Y(n10155) );
  OR2X1_RVT U10041 ( .A1(n12865), .A2(n12263), .Y(n9756) );
  OR2X1_RVT U10042 ( .A1(n9840), .A2(n9890), .Y(n10154) );
  OR2X1_RVT U10043 ( .A1(n12853), .A2(n10156), .Y(n9890) );
  OR2X1_RVT U10044 ( .A1(n10157), .A2(n12246), .Y(n10150) );
  AND4X1_RVT U10045 ( .A1(n10158), .A2(n10159), .A3(n10160), .A4(n10161), .Y(
        n10157) );
  OR2X1_RVT U10046 ( .A1(n10015), .A2(n9788), .Y(n10160) );
  OR2X1_RVT U10047 ( .A1(n10162), .A2(n9785), .Y(n10159) );
  OR2X1_RVT U10048 ( .A1(n12862), .A2(n9740), .Y(n10158) );
  OR2X1_RVT U10049 ( .A1(n10163), .A2(n12247), .Y(n10149) );
  AND2X1_RVT U10050 ( .A1(n10164), .A2(n10165), .Y(n10163) );
  OR2X1_RVT U10051 ( .A1(n10015), .A2(n9740), .Y(n10165) );
  AND2X1_RVT U10052 ( .A1(n10166), .A2(n10016), .Y(n10164) );
  OR2X1_RVT U10053 ( .A1(n9788), .A2(n10167), .Y(n10016) );
  OR2X1_RVT U10054 ( .A1(n12853), .A2(n12865), .Y(n10167) );
  OR2X1_RVT U10055 ( .A1(n10168), .A2(n12254), .Y(n10148) );
  AND4X1_RVT U10056 ( .A1(n10169), .A2(n10003), .A3(n9812), .A4(n9784), .Y(
        n10168) );
  OR2X1_RVT U10057 ( .A1(n9809), .A2(n10170), .Y(n9784) );
  OR2X1_RVT U10058 ( .A1(n12855), .A2(n9746), .Y(n10170) );
  OR2X1_RVT U10059 ( .A1(n9871), .A2(n9905), .Y(n9812) );
  OR2X1_RVT U10060 ( .A1(n9790), .A2(n10171), .Y(n10003) );
  OR2X1_RVT U10061 ( .A1(n12278), .A2(n12247), .Y(n10171) );
  OR2X1_RVT U10062 ( .A1(n9749), .A2(n10172), .Y(n10169) );
  OR2X1_RVT U10063 ( .A1(n10173), .A2(n12252), .Y(n10172) );
  AND4X1_RVT U10064 ( .A1(n10174), .A2(n10175), .A3(n10176), .A4(n10177), .Y(
        n10097) );
  AND2X1_RVT U10065 ( .A1(n10178), .A2(n10179), .Y(n10177) );
  AND2X1_RVT U10066 ( .A1(n10180), .A2(n10181), .Y(n10178) );
  OR2X1_RVT U10067 ( .A1(n9781), .A2(n10135), .Y(n10181) );
  OR2X1_RVT U10068 ( .A1(n9793), .A2(n10182), .Y(n10135) );
  OR2X1_RVT U10069 ( .A1(n12854), .A2(n12856), .Y(n10182) );
  OR2X1_RVT U10070 ( .A1(n12861), .A2(n10183), .Y(n10180) );
  OR2X1_RVT U10071 ( .A1(n12263), .A2(n10184), .Y(n10176) );
  OR2X1_RVT U10072 ( .A1(n12864), .A2(n10185), .Y(n10175) );
  OR2X1_RVT U10073 ( .A1(n9793), .A2(n10186), .Y(n10174) );
  AND4X1_RVT U10074 ( .A1(n10188), .A2(n10189), .A3(n10190), .A4(n10191), .Y(
        n10187) );
  AND4X1_RVT U10075 ( .A1(n10192), .A2(n10193), .A3(n10194), .A4(n10195), .Y(
        n10191) );
  AND4X1_RVT U10076 ( .A1(n10196), .A2(n10197), .A3(n9710), .A4(n10198), .Y(
        n10195) );
  OR2X1_RVT U10077 ( .A1(n9851), .A2(n10199), .Y(n9710) );
  OR2X1_RVT U10078 ( .A1(n9942), .A2(n96), .Y(n10199) );
  OR2X1_RVT U10079 ( .A1(n9714), .A2(n10200), .Y(n10197) );
  OR2X1_RVT U10080 ( .A1(n12859), .A2(n12862), .Y(n10200) );
  OR2X1_RVT U10081 ( .A1(n9977), .A2(n10201), .Y(n10196) );
  OR2X1_RVT U10082 ( .A1(n10202), .A2(n9751), .Y(n10201) );
  AND2X1_RVT U10083 ( .A1(n12267), .A2(n9851), .Y(n10202) );
  OR2X1_RVT U10084 ( .A1(n10203), .A2(n12273), .Y(n10194) );
  AND2X1_RVT U10085 ( .A1(n9992), .A2(n10143), .Y(n10203) );
  OR2X1_RVT U10086 ( .A1(n96), .A2(n10204), .Y(n10143) );
  OR2X1_RVT U10087 ( .A1(n12246), .A2(n12858), .Y(n10204) );
  OR2X1_RVT U10088 ( .A1(n9781), .A2(n10205), .Y(n9992) );
  OR2X1_RVT U10089 ( .A1(n12856), .A2(n9773), .Y(n10205) );
  OR2X1_RVT U10090 ( .A1(n10206), .A2(n9731), .Y(n10193) );
  AND2X1_RVT U10091 ( .A1(n10207), .A2(n9936), .Y(n10206) );
  OR2X1_RVT U10092 ( .A1(n9837), .A2(n9831), .Y(n10192) );
  AND4X1_RVT U10093 ( .A1(n10208), .A2(n10209), .A3(n10210), .A4(n10211), .Y(
        n10190) );
  AND2X1_RVT U10094 ( .A1(n10212), .A2(n10213), .Y(n10211) );
  OR2X1_RVT U10095 ( .A1(n10214), .A2(n12267), .Y(n10213) );
  AND2X1_RVT U10096 ( .A1(n10215), .A2(n9804), .Y(n10214) );
  AND2X1_RVT U10097 ( .A1(n10216), .A2(n10217), .Y(n10212) );
  OR2X1_RVT U10098 ( .A1(n10218), .A2(n9787), .Y(n10217) );
  AND2X1_RVT U10099 ( .A1(n9758), .A2(n9730), .Y(n10218) );
  OR2X1_RVT U10100 ( .A1(n12864), .A2(n9829), .Y(n9758) );
  OR2X1_RVT U10101 ( .A1(n10219), .A2(n9840), .Y(n10216) );
  AND2X1_RVT U10102 ( .A1(n10111), .A2(n10220), .Y(n10219) );
  OR2X1_RVT U10103 ( .A1(n12865), .A2(n9868), .Y(n10111) );
  OR2X1_RVT U10104 ( .A1(n10221), .A2(n12856), .Y(n10210) );
  AND2X1_RVT U10105 ( .A1(n9735), .A2(n10222), .Y(n10221) );
  OR2X1_RVT U10106 ( .A1(n9871), .A2(n9795), .Y(n10222) );
  OR2X1_RVT U10107 ( .A1(n9774), .A2(n9977), .Y(n9735) );
  OR2X1_RVT U10108 ( .A1(n10223), .A2(n94), .Y(n10209) );
  AND2X1_RVT U10109 ( .A1(n9785), .A2(n10224), .Y(n10223) );
  OR2X1_RVT U10110 ( .A1(n10225), .A2(n12251), .Y(n10224) );
  AND2X1_RVT U10111 ( .A1(n10226), .A2(n10227), .Y(n10225) );
  OR2X1_RVT U10112 ( .A1(n12857), .A2(n9768), .Y(n10227) );
  OR2X1_RVT U10113 ( .A1(n12278), .A2(n9871), .Y(n9785) );
  OR2X1_RVT U10114 ( .A1(n10228), .A2(n9855), .Y(n10208) );
  AND2X1_RVT U10115 ( .A1(n9788), .A2(n9833), .Y(n10228) );
  OR2X1_RVT U10116 ( .A1(n12853), .A2(n9716), .Y(n9833) );
  AND4X1_RVT U10117 ( .A1(n10229), .A2(n10230), .A3(n10231), .A4(n10232), .Y(
        n10189) );
  AND4X1_RVT U10118 ( .A1(n10233), .A2(n10234), .A3(n10235), .A4(n10236), .Y(
        n10232) );
  OR2X1_RVT U10119 ( .A1(n10237), .A2(n12864), .Y(n10236) );
  AND2X1_RVT U10120 ( .A1(n9891), .A2(n10238), .Y(n10237) );
  OR2X1_RVT U10121 ( .A1(n12275), .A2(n9740), .Y(n10238) );
  OR2X1_RVT U10122 ( .A1(n10239), .A2(n9733), .Y(n10235) );
  AND2X1_RVT U10123 ( .A1(n10240), .A2(n10241), .Y(n10239) );
  OR2X1_RVT U10124 ( .A1(n10242), .A2(n9768), .Y(n10241) );
  AND2X1_RVT U10125 ( .A1(n9793), .A2(n9781), .Y(n10242) );
  AND2X1_RVT U10126 ( .A1(n9795), .A2(n10116), .Y(n10240) );
  OR2X1_RVT U10127 ( .A1(n12276), .A2(n9933), .Y(n10116) );
  OR2X1_RVT U10128 ( .A1(n10243), .A2(n12265), .Y(n10234) );
  AND2X1_RVT U10129 ( .A1(n10244), .A2(n10245), .Y(n10243) );
  OR2X1_RVT U10130 ( .A1(n9781), .A2(n10246), .Y(n10245) );
  AND2X1_RVT U10131 ( .A1(n9863), .A2(n10136), .Y(n10244) );
  OR2X1_RVT U10132 ( .A1(n9773), .A2(n9948), .Y(n10136) );
  OR2X1_RVT U10133 ( .A1(n9746), .A2(n10247), .Y(n9863) );
  OR2X1_RVT U10134 ( .A1(n10248), .A2(n9716), .Y(n10233) );
  AND4X1_RVT U10135 ( .A1(n10249), .A2(n10250), .A3(n10251), .A4(n10184), .Y(
        n10248) );
  OR2X1_RVT U10136 ( .A1(n9809), .A2(n10252), .Y(n10184) );
  OR2X1_RVT U10137 ( .A1(n12246), .A2(n9773), .Y(n10252) );
  OR2X1_RVT U10138 ( .A1(n12861), .A2(n10015), .Y(n10250) );
  OR2X1_RVT U10139 ( .A1(n9774), .A2(n9871), .Y(n10249) );
  OR2X1_RVT U10140 ( .A1(n9942), .A2(n9984), .Y(n10231) );
  OR2X1_RVT U10141 ( .A1(n10253), .A2(n12249), .Y(n10230) );
  AND4X1_RVT U10142 ( .A1(n10254), .A2(n10255), .A3(n9818), .A4(n9916), .Y(
        n10253) );
  OR2X1_RVT U10143 ( .A1(n9740), .A2(n9905), .Y(n9916) );
  OR2X1_RVT U10144 ( .A1(n12861), .A2(n94), .Y(n9905) );
  OR2X1_RVT U10145 ( .A1(n9733), .A2(n9797), .Y(n9818) );
  OR2X1_RVT U10146 ( .A1(n12853), .A2(n10247), .Y(n10229) );
  AND4X1_RVT U10147 ( .A1(n10256), .A2(n10257), .A3(n10258), .A4(n10259), .Y(
        n10188) );
  OR2X1_RVT U10148 ( .A1(n12254), .A2(n10260), .Y(n10259) );
  AND2X1_RVT U10149 ( .A1(n10261), .A2(n10262), .Y(n10258) );
  OR2X1_RVT U10150 ( .A1(n12275), .A2(n9936), .Y(n10262) );
  OR2X1_RVT U10151 ( .A1(n9723), .A2(n9797), .Y(n10261) );
  OR2X1_RVT U10152 ( .A1(n96), .A2(n9754), .Y(n9797) );
  OR2X1_RVT U10153 ( .A1(n12278), .A2(n9915), .Y(n10257) );
  OR2X1_RVT U10154 ( .A1(n9790), .A2(n10263), .Y(n9915) );
  AND2X1_RVT U10155 ( .A1(n10264), .A2(n10265), .Y(n10256) );
  OR2X1_RVT U10156 ( .A1(n12247), .A2(n10266), .Y(n10265) );
  OR2X1_RVT U10157 ( .A1(n9793), .A2(n9742), .Y(n10264) );
  OR2X1_RVT U10158 ( .A1(n9716), .A2(n10001), .Y(n9742) );
  AND4X1_RVT U10159 ( .A1(n10268), .A2(n10269), .A3(n10270), .A4(n10271), .Y(
        n10267) );
  AND4X1_RVT U10160 ( .A1(n10272), .A2(n10273), .A3(n10274), .A4(n10275), .Y(
        n10271) );
  AND4X1_RVT U10161 ( .A1(n9929), .A2(n10198), .A3(n10276), .A4(n10277), .Y(
        n10275) );
  OR2X1_RVT U10162 ( .A1(n10278), .A2(n10279), .Y(n10198) );
  OR2X1_RVT U10163 ( .A1(n9714), .A2(n9984), .Y(n9929) );
  OR2X1_RVT U10164 ( .A1(n12862), .A2(n12263), .Y(n9984) );
  AND4X1_RVT U10165 ( .A1(n10266), .A2(n10132), .A3(n10255), .A4(n9711), .Y(
        n10274) );
  OR2X1_RVT U10166 ( .A1(n10280), .A2(n9901), .Y(n9711) );
  OR2X1_RVT U10167 ( .A1(n9716), .A2(n10281), .Y(n10255) );
  OR2X1_RVT U10168 ( .A1(n9749), .A2(n94), .Y(n10132) );
  OR2X1_RVT U10169 ( .A1(n9740), .A2(n10282), .Y(n10266) );
  OR2X1_RVT U10170 ( .A1(n12253), .A2(n12273), .Y(n10282) );
  AND4X1_RVT U10171 ( .A1(n10283), .A2(n10284), .A3(n10285), .A4(n10286), .Y(
        n10273) );
  OR2X1_RVT U10172 ( .A1(n9993), .A2(n10287), .Y(n10286) );
  OR2X1_RVT U10173 ( .A1(n12273), .A2(n9773), .Y(n10287) );
  OR2X1_RVT U10174 ( .A1(n9902), .A2(n10288), .Y(n10285) );
  OR2X1_RVT U10175 ( .A1(n12863), .A2(n9790), .Y(n10288) );
  OR2X1_RVT U10176 ( .A1(n10207), .A2(n10289), .Y(n10284) );
  OR2X1_RVT U10177 ( .A1(n10290), .A2(n9787), .Y(n10289) );
  OR2X1_RVT U10178 ( .A1(n12270), .A2(n10291), .Y(n10283) );
  OR2X1_RVT U10179 ( .A1(n10292), .A2(n12253), .Y(n10291) );
  AND2X1_RVT U10180 ( .A1(n10001), .A2(n10293), .Y(n10292) );
  AND2X1_RVT U10181 ( .A1(n10294), .A2(n10295), .Y(n10272) );
  OR2X1_RVT U10182 ( .A1(n10296), .A2(n9768), .Y(n10295) );
  AND2X1_RVT U10183 ( .A1(n10297), .A2(n10298), .Y(n10296) );
  OR2X1_RVT U10184 ( .A1(n12252), .A2(n9961), .Y(n10298) );
  OR2X1_RVT U10185 ( .A1(n12256), .A2(n10115), .Y(n10297) );
  AND2X1_RVT U10186 ( .A1(n10299), .A2(n10300), .Y(n10294) );
  OR2X1_RVT U10187 ( .A1(n10301), .A2(n9807), .Y(n10300) );
  AND2X1_RVT U10188 ( .A1(n10302), .A2(n10303), .Y(n10301) );
  OR2X1_RVT U10189 ( .A1(n12259), .A2(n104), .Y(n10303) );
  NAND2X1_RVT U10190 ( .A1(n9790), .A2(n12855), .Y(n10302) );
  OR2X1_RVT U10191 ( .A1(n10304), .A2(n96), .Y(n10299) );
  AND2X1_RVT U10192 ( .A1(n10014), .A2(n9891), .Y(n10304) );
  OR2X1_RVT U10193 ( .A1(n9740), .A2(n10305), .Y(n9891) );
  OR2X1_RVT U10194 ( .A1(n12866), .A2(n12248), .Y(n10305) );
  AND4X1_RVT U10195 ( .A1(n9908), .A2(n10306), .A3(n10179), .A4(n10307), .Y(
        n10270) );
  AND4X1_RVT U10196 ( .A1(n10308), .A2(n10309), .A3(n10310), .A4(n10311), .Y(
        n10307) );
  OR2X1_RVT U10197 ( .A1(n9871), .A2(n9792), .Y(n10311) );
  OR2X1_RVT U10198 ( .A1(n9809), .A2(n9838), .Y(n10310) );
  OR2X1_RVT U10199 ( .A1(n12854), .A2(n10142), .Y(n10309) );
  OR2X1_RVT U10200 ( .A1(n9787), .A2(n9769), .Y(n10142) );
  OR2X1_RVT U10201 ( .A1(n12862), .A2(n9851), .Y(n9769) );
  OR2X1_RVT U10202 ( .A1(n12262), .A2(n9892), .Y(n10308) );
  OR2X1_RVT U10203 ( .A1(n9773), .A2(n10001), .Y(n9892) );
  OR2X1_RVT U10204 ( .A1(n12246), .A2(n9977), .Y(n10001) );
  AND2X1_RVT U10205 ( .A1(n10312), .A2(n10313), .Y(n10179) );
  OR2X1_RVT U10206 ( .A1(n10314), .A2(n9840), .Y(n10313) );
  OR2X1_RVT U10207 ( .A1(n12272), .A2(n96), .Y(n10314) );
  OR2X1_RVT U10208 ( .A1(n10315), .A2(n9723), .Y(n10312) );
  OR2X1_RVT U10209 ( .A1(n12853), .A2(n9840), .Y(n9723) );
  OR2X1_RVT U10210 ( .A1(n9737), .A2(n9787), .Y(n10315) );
  OR2X1_RVT U10211 ( .A1(n12254), .A2(n10185), .Y(n10306) );
  AND2X1_RVT U10212 ( .A1(n10316), .A2(n10317), .Y(n9908) );
  OR2X1_RVT U10213 ( .A1(n9791), .A2(n9829), .Y(n10317) );
  OR2X1_RVT U10214 ( .A1(n10318), .A2(n10319), .Y(n10316) );
  AND4X1_RVT U10215 ( .A1(n10320), .A2(n10321), .A3(n10322), .A4(n10323), .Y(
        n10269) );
  OR2X1_RVT U10216 ( .A1(n10324), .A2(n9977), .Y(n10323) );
  AND2X1_RVT U10217 ( .A1(n10325), .A2(n9986), .Y(n10324) );
  OR2X1_RVT U10218 ( .A1(n12260), .A2(n10281), .Y(n9986) );
  OR2X1_RVT U10219 ( .A1(n10326), .A2(n12859), .Y(n10322) );
  AND2X1_RVT U10220 ( .A1(n9914), .A2(n9879), .Y(n10326) );
  OR2X1_RVT U10221 ( .A1(n12853), .A2(n9855), .Y(n9879) );
  OR2X1_RVT U10222 ( .A1(n10327), .A2(n9934), .Y(n10321) );
  AND2X1_RVT U10223 ( .A1(n10328), .A2(n10329), .Y(n10327) );
  OR2X1_RVT U10224 ( .A1(n12249), .A2(n9793), .Y(n10329) );
  AND2X1_RVT U10225 ( .A1(n10330), .A2(n9831), .Y(n10328) );
  OR2X1_RVT U10226 ( .A1(n94), .A2(n9790), .Y(n10330) );
  OR2X1_RVT U10227 ( .A1(n10331), .A2(n9731), .Y(n10320) );
  AND2X1_RVT U10228 ( .A1(n10332), .A2(n10333), .Y(n10331) );
  NAND2X1_RVT U10229 ( .A1(n9716), .A2(n10173), .Y(n10333) );
  AND2X1_RVT U10230 ( .A1(n10334), .A2(n9944), .Y(n10332) );
  OR2X1_RVT U10231 ( .A1(n9877), .A2(n10281), .Y(n9944) );
  OR2X1_RVT U10232 ( .A1(n12269), .A2(n10335), .Y(n10334) );
  AND4X1_RVT U10233 ( .A1(n10336), .A2(n10337), .A3(n10338), .A4(n10339), .Y(
        n10268) );
  OR2X1_RVT U10234 ( .A1(n10340), .A2(n9754), .Y(n10339) );
  AND2X1_RVT U10235 ( .A1(n10341), .A2(n9895), .Y(n10340) );
  AND2X1_RVT U10236 ( .A1(n10342), .A2(n9917), .Y(n10341) );
  OR2X1_RVT U10237 ( .A1(n96), .A2(n10319), .Y(n9917) );
  OR2X1_RVT U10238 ( .A1(n12248), .A2(n9851), .Y(n10319) );
  OR2X1_RVT U10239 ( .A1(n10343), .A2(n12265), .Y(n10338) );
  AND2X1_RVT U10240 ( .A1(n10344), .A2(n10345), .Y(n10343) );
  OR2X1_RVT U10241 ( .A1(n10346), .A2(n12851), .Y(n10345) );
  AND2X1_RVT U10242 ( .A1(n10347), .A2(n10348), .Y(n10346) );
  OR2X1_RVT U10243 ( .A1(n12247), .A2(n10207), .Y(n10348) );
  OR2X1_RVT U10244 ( .A1(n12858), .A2(n9774), .Y(n10347) );
  AND2X1_RVT U10245 ( .A1(n10349), .A2(n10350), .Y(n10344) );
  OR2X1_RVT U10246 ( .A1(n9740), .A2(n10351), .Y(n10349) );
  OR2X1_RVT U10247 ( .A1(n10352), .A2(n9774), .Y(n10337) );
  AND4X1_RVT U10248 ( .A1(n10353), .A2(n10354), .A3(n10355), .A4(n9740), .Y(
        n10352) );
  OR2X1_RVT U10249 ( .A1(n12859), .A2(n9790), .Y(n10355) );
  OR2X1_RVT U10250 ( .A1(n12259), .A2(n9809), .Y(n10354) );
  OR2X1_RVT U10251 ( .A1(n9862), .A2(n9840), .Y(n10353) );
  OR2X1_RVT U10252 ( .A1(n10356), .A2(n9716), .Y(n10336) );
  AND4X1_RVT U10253 ( .A1(n10220), .A2(n10357), .A3(n9939), .A4(n9855), .Y(
        n10356) );
  OR2X1_RVT U10254 ( .A1(n9809), .A2(n10351), .Y(n9939) );
  OR2X1_RVT U10255 ( .A1(n9977), .A2(n10263), .Y(n10357) );
  OR2X1_RVT U10256 ( .A1(n12253), .A2(n9942), .Y(n10220) );
  AND4X1_RVT U10257 ( .A1(n10359), .A2(n10360), .A3(n10361), .A4(n10362), .Y(
        n10358) );
  AND4X1_RVT U10258 ( .A1(n9792), .A2(n10107), .A3(n10363), .A4(n10364), .Y(
        n10362) );
  AND4X1_RVT U10259 ( .A1(n10186), .A2(n10131), .A3(n10276), .A4(n10277), .Y(
        n10364) );
  OR2X1_RVT U10260 ( .A1(n10279), .A2(n9713), .Y(n10277) );
  OR2X1_RVT U10261 ( .A1(n12857), .A2(n9831), .Y(n9713) );
  OR2X1_RVT U10262 ( .A1(n9730), .A2(n10318), .Y(n10276) );
  OR2X1_RVT U10263 ( .A1(n12862), .A2(n12267), .Y(n10318) );
  OR2X1_RVT U10264 ( .A1(n12851), .A2(n9851), .Y(n9730) );
  OR2X1_RVT U10265 ( .A1(n12863), .A2(n9749), .Y(n10131) );
  OR2X1_RVT U10266 ( .A1(n12276), .A2(n12260), .Y(n9749) );
  OR2X1_RVT U10267 ( .A1(n9871), .A2(n10365), .Y(n10186) );
  OR2X1_RVT U10268 ( .A1(n12267), .A2(n9775), .Y(n10365) );
  OR2X1_RVT U10269 ( .A1(n9773), .A2(n10366), .Y(n10363) );
  OR2X1_RVT U10270 ( .A1(n9901), .A2(n12258), .Y(n10366) );
  OR2X1_RVT U10271 ( .A1(n9840), .A2(n10367), .Y(n10107) );
  OR2X1_RVT U10272 ( .A1(n9774), .A2(n12265), .Y(n10367) );
  OR2X1_RVT U10273 ( .A1(n12855), .A2(n10278), .Y(n9792) );
  OR2X1_RVT U10274 ( .A1(n12260), .A2(n9791), .Y(n10278) );
  AND4X1_RVT U10275 ( .A1(n10368), .A2(n10369), .A3(n10370), .A4(n10371), .Y(
        n10361) );
  AND4X1_RVT U10276 ( .A1(n10372), .A2(n10373), .A3(n10374), .A4(n10375), .Y(
        n10371) );
  OR2X1_RVT U10277 ( .A1(n9807), .A2(n10376), .Y(n10375) );
  OR2X1_RVT U10278 ( .A1(n12249), .A2(n9877), .Y(n10376) );
  OR2X1_RVT U10279 ( .A1(n9790), .A2(n10377), .Y(n10374) );
  OR2X1_RVT U10280 ( .A1(n10378), .A2(n9754), .Y(n10377) );
  AND2X1_RVT U10281 ( .A1(n9733), .A2(n9793), .Y(n10378) );
  OR2X1_RVT U10282 ( .A1(n10379), .A2(n10380), .Y(n10373) );
  AND2X1_RVT U10283 ( .A1(n9948), .A2(n9904), .Y(n10379) );
  OR2X1_RVT U10284 ( .A1(n12856), .A2(n104), .Y(n9904) );
  OR2X1_RVT U10285 ( .A1(n12852), .A2(n12270), .Y(n9948) );
  OR2X1_RVT U10286 ( .A1(n10381), .A2(n9788), .Y(n10372) );
  AND2X1_RVT U10287 ( .A1(n10263), .A2(n10382), .Y(n10381) );
  OR2X1_RVT U10288 ( .A1(n12854), .A2(n96), .Y(n10382) );
  OR2X1_RVT U10289 ( .A1(n10383), .A2(n12272), .Y(n10370) );
  AND2X1_RVT U10290 ( .A1(n10254), .A2(n10384), .Y(n10383) );
  OR2X1_RVT U10291 ( .A1(n9781), .A2(n10207), .Y(n10384) );
  OR2X1_RVT U10292 ( .A1(n12253), .A2(n9993), .Y(n10254) );
  OR2X1_RVT U10293 ( .A1(n12858), .A2(n9781), .Y(n9993) );
  OR2X1_RVT U10294 ( .A1(n10385), .A2(n9942), .Y(n10369) );
  AND2X1_RVT U10295 ( .A1(n9895), .A2(n10246), .Y(n10385) );
  OR2X1_RVT U10296 ( .A1(n9751), .A2(n9840), .Y(n9895) );
  OR2X1_RVT U10297 ( .A1(n10386), .A2(n9831), .Y(n10368) );
  AND2X1_RVT U10298 ( .A1(n9794), .A2(n9796), .Y(n10386) );
  AND4X1_RVT U10299 ( .A1(n10387), .A2(n10388), .A3(n10389), .A4(n10390), .Y(
        n10360) );
  AND4X1_RVT U10300 ( .A1(n10391), .A2(n10392), .A3(n10393), .A4(n10394), .Y(
        n10390) );
  OR2X1_RVT U10301 ( .A1(n10395), .A2(n12256), .Y(n10394) );
  AND2X1_RVT U10302 ( .A1(n9722), .A2(n10014), .Y(n10395) );
  OR2X1_RVT U10303 ( .A1(n9871), .A2(n9902), .Y(n10014) );
  OR2X1_RVT U10304 ( .A1(n12259), .A2(n9754), .Y(n9902) );
  OR2X1_RVT U10305 ( .A1(n12263), .A2(n10396), .Y(n9722) );
  OR2X1_RVT U10306 ( .A1(n12246), .A2(n12252), .Y(n10396) );
  OR2X1_RVT U10307 ( .A1(n10397), .A2(n12270), .Y(n10393) );
  AND2X1_RVT U10308 ( .A1(n10110), .A2(n10398), .Y(n10397) );
  OR2X1_RVT U10309 ( .A1(n12275), .A2(n94), .Y(n10398) );
  OR2X1_RVT U10310 ( .A1(n12273), .A2(n9838), .Y(n10110) );
  OR2X1_RVT U10311 ( .A1(n10399), .A2(n12251), .Y(n10392) );
  AND2X1_RVT U10312 ( .A1(n10128), .A2(n10400), .Y(n10399) );
  OR2X1_RVT U10313 ( .A1(n12276), .A2(n9774), .Y(n10400) );
  OR2X1_RVT U10314 ( .A1(n9716), .A2(n10401), .Y(n10128) );
  OR2X1_RVT U10315 ( .A1(n10402), .A2(n9775), .Y(n10391) );
  AND2X1_RVT U10316 ( .A1(n10403), .A2(n10404), .Y(n10402) );
  OR2X1_RVT U10317 ( .A1(n9831), .A2(n12273), .Y(n10404) );
  AND2X1_RVT U10318 ( .A1(n10405), .A2(n9807), .Y(n10403) );
  OR2X1_RVT U10319 ( .A1(n9793), .A2(n9754), .Y(n9807) );
  OR2X1_RVT U10320 ( .A1(n12248), .A2(n9838), .Y(n10405) );
  OR2X1_RVT U10321 ( .A1(n12866), .A2(n9793), .Y(n9838) );
  OR2X1_RVT U10322 ( .A1(n10406), .A2(n9851), .Y(n10389) );
  AND4X1_RVT U10323 ( .A1(n10407), .A2(n10408), .A3(n10004), .A4(n9914), .Y(
        n10406) );
  OR2X1_RVT U10324 ( .A1(n9977), .A2(n10156), .Y(n9914) );
  OR2X1_RVT U10325 ( .A1(n9809), .A2(n10335), .Y(n10004) );
  OR2X1_RVT U10326 ( .A1(n12254), .A2(n12247), .Y(n10335) );
  OR2X1_RVT U10327 ( .A1(n96), .A2(n9731), .Y(n10408) );
  OR2X1_RVT U10328 ( .A1(n94), .A2(n12273), .Y(n10407) );
  OR2X1_RVT U10329 ( .A1(n10409), .A2(n9787), .Y(n10388) );
  AND2X1_RVT U10330 ( .A1(n10410), .A2(n9808), .Y(n10409) );
  AND2X1_RVT U10331 ( .A1(n10342), .A2(n10137), .Y(n10410) );
  OR2X1_RVT U10332 ( .A1(n10411), .A2(n12863), .Y(n10137) );
  AND2X1_RVT U10333 ( .A1(n9829), .A2(n10412), .Y(n10411) );
  OR2X1_RVT U10334 ( .A1(n12251), .A2(n9716), .Y(n10412) );
  OR2X1_RVT U10335 ( .A1(n9877), .A2(n10015), .Y(n10342) );
  OR2X1_RVT U10336 ( .A1(n9862), .A2(n9751), .Y(n10015) );
  OR2X1_RVT U10337 ( .A1(n10413), .A2(n9855), .Y(n10387) );
  AND2X1_RVT U10338 ( .A1(n10414), .A2(n12259), .Y(n10413) );
  AND2X1_RVT U10339 ( .A1(n10415), .A2(n10115), .Y(n10414) );
  OR2X1_RVT U10340 ( .A1(n9877), .A2(n9977), .Y(n10415) );
  AND4X1_RVT U10341 ( .A1(n10416), .A2(n10417), .A3(n10418), .A4(n10419), .Y(
        n10359) );
  AND2X1_RVT U10342 ( .A1(n10420), .A2(n10421), .Y(n10419) );
  OR2X1_RVT U10343 ( .A1(n12859), .A2(n9957), .Y(n10421) );
  OR2X1_RVT U10344 ( .A1(n12267), .A2(n10422), .Y(n9957) );
  OR2X1_RVT U10345 ( .A1(n9773), .A2(n9862), .Y(n10422) );
  AND2X1_RVT U10346 ( .A1(n10423), .A2(n10424), .Y(n10420) );
  OR2X1_RVT U10347 ( .A1(n9746), .A2(n9757), .Y(n10424) );
  OR2X1_RVT U10348 ( .A1(n9790), .A2(n9985), .Y(n9757) );
  OR2X1_RVT U10349 ( .A1(n12855), .A2(n9751), .Y(n9985) );
  OR2X1_RVT U10350 ( .A1(n9793), .A2(n9870), .Y(n10423) );
  OR2X1_RVT U10351 ( .A1(n9781), .A2(n10425), .Y(n9870) );
  OR2X1_RVT U10352 ( .A1(n9781), .A2(n9961), .Y(n10418) );
  OR2X1_RVT U10353 ( .A1(n96), .A2(n12269), .Y(n9961) );
  OR2X1_RVT U10354 ( .A1(n10426), .A2(n9737), .Y(n10417) );
  AND4X1_RVT U10355 ( .A1(n10427), .A2(n10428), .A3(n10429), .A4(n10430), .Y(
        n10426) );
  OR2X1_RVT U10356 ( .A1(n12853), .A2(n10431), .Y(n10429) );
  OR2X1_RVT U10357 ( .A1(n10432), .A2(n12860), .Y(n10431) );
  AND2X1_RVT U10358 ( .A1(n9788), .A2(n10433), .Y(n10432) );
  OR2X1_RVT U10359 ( .A1(n12262), .A2(n10434), .Y(n10428) );
  OR2X1_RVT U10360 ( .A1(n10173), .A2(n9731), .Y(n10434) );
  OR2X1_RVT U10361 ( .A1(n9714), .A2(n9740), .Y(n10427) );
  OR2X1_RVT U10362 ( .A1(n12857), .A2(n9840), .Y(n9740) );
  OR2X1_RVT U10363 ( .A1(n10293), .A2(n10207), .Y(n10416) );
  OR2X1_RVT U10364 ( .A1(n12278), .A2(n9751), .Y(n10207) );
  AND4X1_RVT U10365 ( .A1(n10436), .A2(n10437), .A3(n10438), .A4(n10439), .Y(
        n10435) );
  AND4X1_RVT U10366 ( .A1(n10440), .A2(n10441), .A3(n10442), .A4(n10443), .Y(
        n10439) );
  AND4X1_RVT U10367 ( .A1(n10444), .A2(n10445), .A3(n10446), .A4(n10447), .Y(
        n10443) );
  OR2X1_RVT U10368 ( .A1(n10281), .A2(n10425), .Y(n10447) );
  OR2X1_RVT U10369 ( .A1(n12856), .A2(n12272), .Y(n10425) );
  OR2X1_RVT U10370 ( .A1(n12246), .A2(n12256), .Y(n10281) );
  OR2X1_RVT U10371 ( .A1(n10448), .A2(n9788), .Y(n10446) );
  AND2X1_RVT U10372 ( .A1(n9734), .A2(n10380), .Y(n10448) );
  OR2X1_RVT U10373 ( .A1(n96), .A2(n10449), .Y(n9734) );
  OR2X1_RVT U10374 ( .A1(n12246), .A2(n12853), .Y(n10449) );
  OR2X1_RVT U10375 ( .A1(n10450), .A2(n9716), .Y(n10445) );
  OR2X1_RVT U10376 ( .A1(n12260), .A2(n9877), .Y(n9716) );
  AND2X1_RVT U10377 ( .A1(n9852), .A2(n10451), .Y(n10450) );
  OR2X1_RVT U10378 ( .A1(n9731), .A2(n9933), .Y(n10451) );
  OR2X1_RVT U10379 ( .A1(n12264), .A2(n12252), .Y(n9731) );
  OR2X1_RVT U10380 ( .A1(n9977), .A2(n10452), .Y(n9852) );
  OR2X1_RVT U10381 ( .A1(n12864), .A2(n12267), .Y(n10452) );
  OR2X1_RVT U10382 ( .A1(n10453), .A2(n9775), .Y(n10444) );
  AND2X1_RVT U10383 ( .A1(n10251), .A2(n10454), .Y(n10453) );
  OR2X1_RVT U10384 ( .A1(n10455), .A2(n12853), .Y(n10454) );
  AND2X1_RVT U10385 ( .A1(n9831), .A2(n10263), .Y(n10455) );
  OR2X1_RVT U10386 ( .A1(n12861), .A2(n9793), .Y(n10263) );
  OR2X1_RVT U10387 ( .A1(n12273), .A2(n10456), .Y(n10251) );
  OR2X1_RVT U10388 ( .A1(n12866), .A2(n12862), .Y(n10456) );
  OR2X1_RVT U10389 ( .A1(n10457), .A2(n12251), .Y(n10442) );
  AND2X1_RVT U10390 ( .A1(n10458), .A2(n10459), .Y(n10457) );
  OR2X1_RVT U10391 ( .A1(n10460), .A2(n9877), .Y(n10459) );
  AND2X1_RVT U10392 ( .A1(n9942), .A2(n10461), .Y(n10460) );
  OR2X1_RVT U10393 ( .A1(n9733), .A2(n9855), .Y(n10458) );
  OR2X1_RVT U10394 ( .A1(n12265), .A2(n9791), .Y(n9855) );
  OR2X1_RVT U10395 ( .A1(n10462), .A2(n12862), .Y(n10441) );
  AND2X1_RVT U10396 ( .A1(n9947), .A2(n10185), .Y(n10462) );
  OR2X1_RVT U10397 ( .A1(n12263), .A2(n10463), .Y(n10185) );
  OR2X1_RVT U10398 ( .A1(n9787), .A2(n12252), .Y(n10463) );
  OR2X1_RVT U10399 ( .A1(n9733), .A2(n10293), .Y(n9947) );
  OR2X1_RVT U10400 ( .A1(n12252), .A2(n12267), .Y(n10293) );
  OR2X1_RVT U10401 ( .A1(n10464), .A2(n12249), .Y(n10440) );
  AND2X1_RVT U10402 ( .A1(n9987), .A2(n10465), .Y(n10464) );
  OR2X1_RVT U10403 ( .A1(n10280), .A2(n9781), .Y(n10465) );
  OR2X1_RVT U10404 ( .A1(n9840), .A2(n10401), .Y(n9987) );
  OR2X1_RVT U10405 ( .A1(n12861), .A2(n96), .Y(n10401) );
  AND2X1_RVT U10406 ( .A1(n12253), .A2(n12864), .Y(n10162) );
  AND4X1_RVT U10407 ( .A1(n10466), .A2(n10467), .A3(n10468), .A4(n10469), .Y(
        n10438) );
  AND4X1_RVT U10408 ( .A1(n10470), .A2(n10471), .A3(n10472), .A4(n10473), .Y(
        n10469) );
  OR2X1_RVT U10409 ( .A1(n10474), .A2(n12258), .Y(n10473) );
  AND2X1_RVT U10410 ( .A1(n9974), .A2(n10124), .Y(n10474) );
  OR2X1_RVT U10411 ( .A1(n9790), .A2(n10380), .Y(n10124) );
  OR2X1_RVT U10412 ( .A1(n12864), .A2(n9787), .Y(n10380) );
  OR2X1_RVT U10413 ( .A1(n12851), .A2(n12248), .Y(n9790) );
  OR2X1_RVT U10414 ( .A1(n12249), .A2(n10156), .Y(n9974) );
  OR2X1_RVT U10415 ( .A1(n12253), .A2(n12267), .Y(n10156) );
  OR2X1_RVT U10416 ( .A1(n10475), .A2(n12860), .Y(n10472) );
  AND2X1_RVT U10417 ( .A1(n10215), .A2(n10476), .Y(n10475) );
  OR2X1_RVT U10418 ( .A1(n10173), .A2(n9804), .Y(n10476) );
  OR2X1_RVT U10419 ( .A1(n9977), .A2(n10477), .Y(n9804) );
  OR2X1_RVT U10420 ( .A1(n12278), .A2(n12254), .Y(n10477) );
  OR2X1_RVT U10421 ( .A1(n12262), .A2(n10478), .Y(n10215) );
  OR2X1_RVT U10422 ( .A1(n9977), .A2(n9773), .Y(n10478) );
  OR2X1_RVT U10423 ( .A1(n10479), .A2(n12866), .Y(n10471) );
  AND2X1_RVT U10424 ( .A1(n10161), .A2(n10011), .Y(n10479) );
  OR2X1_RVT U10425 ( .A1(n9793), .A2(n9829), .Y(n10011) );
  OR2X1_RVT U10426 ( .A1(n12858), .A2(n9977), .Y(n9829) );
  OR2X1_RVT U10427 ( .A1(n10280), .A2(n9809), .Y(n10161) );
  OR2X1_RVT U10428 ( .A1(n12259), .A2(n12863), .Y(n10280) );
  OR2X1_RVT U10429 ( .A1(n10480), .A2(n9851), .Y(n10470) );
  AND2X1_RVT U10430 ( .A1(n10481), .A2(n10482), .Y(n10480) );
  OR2X1_RVT U10431 ( .A1(n9773), .A2(n10279), .Y(n10482) );
  OR2X1_RVT U10432 ( .A1(n12860), .A2(n104), .Y(n10279) );
  AND2X1_RVT U10433 ( .A1(n10483), .A2(n10147), .Y(n10481) );
  OR2X1_RVT U10434 ( .A1(n9781), .A2(n10484), .Y(n10147) );
  OR2X1_RVT U10435 ( .A1(n12275), .A2(n12254), .Y(n10484) );
  OR2X1_RVT U10436 ( .A1(n9837), .A2(n9774), .Y(n10468) );
  OR2X1_RVT U10437 ( .A1(n12853), .A2(n9733), .Y(n9837) );
  OR2X1_RVT U10438 ( .A1(n10485), .A2(n9737), .Y(n10467) );
  AND2X1_RVT U10439 ( .A1(n10486), .A2(n9918), .Y(n10485) );
  AND2X1_RVT U10440 ( .A1(n10487), .A2(n10488), .Y(n9918) );
  OR2X1_RVT U10441 ( .A1(n12263), .A2(n9942), .Y(n10488) );
  OR2X1_RVT U10442 ( .A1(n9840), .A2(n9714), .Y(n10487) );
  OR2X1_RVT U10443 ( .A1(n12248), .A2(n9787), .Y(n9714) );
  AND2X1_RVT U10444 ( .A1(n10489), .A2(n10183), .Y(n10486) );
  OR2X1_RVT U10445 ( .A1(n9871), .A2(n10433), .Y(n10183) );
  OR2X1_RVT U10446 ( .A1(n12855), .A2(n94), .Y(n10433) );
  OR2X1_RVT U10447 ( .A1(n9733), .A2(n9900), .Y(n10489) );
  OR2X1_RVT U10448 ( .A1(n12247), .A2(n10490), .Y(n9900) );
  OR2X1_RVT U10449 ( .A1(n12851), .A2(n12276), .Y(n10490) );
  OR2X1_RVT U10450 ( .A1(n10491), .A2(n12851), .Y(n10466) );
  AND4X1_RVT U10451 ( .A1(n10492), .A2(n10493), .A3(n10494), .A4(n10325), .Y(
        n10491) );
  OR2X1_RVT U10452 ( .A1(n9787), .A2(n10246), .Y(n10325) );
  OR2X1_RVT U10453 ( .A1(n12856), .A2(n12862), .Y(n10246) );
  OR2X1_RVT U10454 ( .A1(n9787), .A2(n10495), .Y(n10494) );
  OR2X1_RVT U10455 ( .A1(n12253), .A2(n12258), .Y(n10495) );
  OR2X1_RVT U10456 ( .A1(n12861), .A2(n9746), .Y(n9787) );
  OR2X1_RVT U10457 ( .A1(n10496), .A2(n9868), .Y(n10493) );
  OR2X1_RVT U10458 ( .A1(n12247), .A2(n9712), .Y(n9868) );
  AND2X1_RVT U10459 ( .A1(n9851), .A2(n10497), .Y(n10496) );
  OR2X1_RVT U10460 ( .A1(n12859), .A2(n9751), .Y(n10497) );
  OR2X1_RVT U10461 ( .A1(n12855), .A2(n12258), .Y(n9851) );
  OR2X1_RVT U10462 ( .A1(n12857), .A2(n10461), .Y(n10492) );
  OR2X1_RVT U10463 ( .A1(n12861), .A2(n9791), .Y(n10461) );
  OR2X1_RVT U10464 ( .A1(n9737), .A2(n94), .Y(n9791) );
  AND4X1_RVT U10465 ( .A1(n10498), .A2(n10499), .A3(n10500), .A4(n10501), .Y(
        n10437) );
  AND4X1_RVT U10466 ( .A1(n10502), .A2(n10503), .A3(n10504), .A4(n10505), .Y(
        n10501) );
  OR2X1_RVT U10467 ( .A1(n9809), .A2(n9936), .Y(n10505) );
  OR2X1_RVT U10468 ( .A1(n12260), .A2(n9831), .Y(n9936) );
  OR2X1_RVT U10469 ( .A1(n12264), .A2(n9977), .Y(n9809) );
  OR2X1_RVT U10470 ( .A1(n9796), .A2(n10351), .Y(n10504) );
  OR2X1_RVT U10471 ( .A1(n12865), .A2(n12247), .Y(n10351) );
  OR2X1_RVT U10472 ( .A1(n9862), .A2(n9788), .Y(n9796) );
  OR2X1_RVT U10473 ( .A1(n9781), .A2(n9808), .Y(n10503) );
  OR2X1_RVT U10474 ( .A1(n12256), .A2(n12269), .Y(n9808) );
  OR2X1_RVT U10475 ( .A1(n12246), .A2(n12852), .Y(n9781) );
  OR2X1_RVT U10476 ( .A1(n104), .A2(n10226), .Y(n10502) );
  OR2X1_RVT U10477 ( .A1(n12254), .A2(n9934), .Y(n10226) );
  OR2X1_RVT U10478 ( .A1(n9751), .A2(n10260), .Y(n10500) );
  OR2X1_RVT U10479 ( .A1(n104), .A2(n10506), .Y(n10260) );
  OR2X1_RVT U10480 ( .A1(n12858), .A2(n12267), .Y(n10506) );
  AND2X1_RVT U10481 ( .A1(n12248), .A2(n12251), .Y(n10290) );
  OR2X1_RVT U10482 ( .A1(n9793), .A2(n9741), .Y(n10499) );
  OR2X1_RVT U10483 ( .A1(n12276), .A2(n10507), .Y(n9741) );
  OR2X1_RVT U10484 ( .A1(n12859), .A2(n12851), .Y(n10507) );
  OR2X1_RVT U10485 ( .A1(n12253), .A2(n9773), .Y(n9793) );
  OR2X1_RVT U10486 ( .A1(n9840), .A2(n10483), .Y(n10498) );
  OR2X1_RVT U10487 ( .A1(n12249), .A2(n9795), .Y(n10483) );
  OR2X1_RVT U10488 ( .A1(n12861), .A2(n12862), .Y(n9795) );
  AND4X1_RVT U10489 ( .A1(n10508), .A2(n9906), .A3(n10509), .A4(n10510), .Y(
        n10436) );
  OR2X1_RVT U10490 ( .A1(n12253), .A2(n10430), .Y(n10510) );
  OR2X1_RVT U10491 ( .A1(n12857), .A2(n9901), .Y(n10430) );
  OR2X1_RVT U10492 ( .A1(n12251), .A2(n9942), .Y(n9901) );
  OR2X1_RVT U10493 ( .A1(n12246), .A2(n9768), .Y(n9942) );
  AND2X1_RVT U10494 ( .A1(n10511), .A2(n10512), .Y(n10509) );
  OR2X1_RVT U10495 ( .A1(n12275), .A2(n10350), .Y(n10512) );
  OR2X1_RVT U10496 ( .A1(n9840), .A2(n9933), .Y(n10350) );
  OR2X1_RVT U10497 ( .A1(n12253), .A2(n12247), .Y(n9933) );
  OR2X1_RVT U10498 ( .A1(n12248), .A2(n9729), .Y(n9768) );
  OR2X1_RVT U10499 ( .A1(n12864), .A2(n10002), .Y(n10511) );
  OR2X1_RVT U10500 ( .A1(n12272), .A2(n10115), .Y(n10002) );
  OR2X1_RVT U10501 ( .A1(n12856), .A2(n12851), .Y(n10115) );
  OR2X1_RVT U10502 ( .A1(n12854), .A2(n12264), .Y(n9712) );
  AND2X1_RVT U10503 ( .A1(n10513), .A2(n10514), .Y(n9906) );
  OR2X1_RVT U10504 ( .A1(n9788), .A2(n9774), .Y(n10514) );
  OR2X1_RVT U10505 ( .A1(n12863), .A2(n9746), .Y(n9774) );
  AND2X1_RVT U10506 ( .A1(n9773), .A2(n9737), .Y(n9826) );
  OR2X1_RVT U10507 ( .A1(n12259), .A2(n9840), .Y(n9788) );
  OR2X1_RVT U10508 ( .A1(n12852), .A2(n9877), .Y(n9840) );
  OR2X1_RVT U10509 ( .A1(n10515), .A2(n9831), .Y(n10513) );
  OR2X1_RVT U10510 ( .A1(n12253), .A2(n94), .Y(n9831) );
  AND2X1_RVT U10511 ( .A1(n12865), .A2(n12246), .Y(n10173) );
  OR2X1_RVT U10512 ( .A1(n12252), .A2(n9934), .Y(n10515) );
  OR2X1_RVT U10513 ( .A1(n12861), .A2(n12269), .Y(n9934) );
  AND2X1_RVT U10514 ( .A1(n10516), .A2(n10517), .Y(n10508) );
  OR2X1_RVT U10515 ( .A1(n9754), .A2(n10166), .Y(n10517) );
  OR2X1_RVT U10516 ( .A1(n12254), .A2(n9794), .Y(n10166) );
  OR2X1_RVT U10517 ( .A1(n12269), .A2(n9871), .Y(n9794) );
  OR2X1_RVT U10518 ( .A1(n12249), .A2(n12252), .Y(n9871) );
  OR2X1_RVT U10519 ( .A1(n12858), .A2(n12856), .Y(n9733) );
  OR2X1_RVT U10520 ( .A1(n12866), .A2(n12860), .Y(n9754) );
  XOR2X1_RVT U10521 ( .A1(key[92]), .A2(state[92]), .Y(n9729) );
  OR2X1_RVT U10522 ( .A1(n9746), .A2(n9875), .Y(n10516) );
  OR2X1_RVT U10523 ( .A1(n9977), .A2(n10247), .Y(n9875) );
  OR2X1_RVT U10524 ( .A1(n12256), .A2(n9775), .Y(n10247) );
  OR2X1_RVT U10525 ( .A1(n12859), .A2(n9877), .Y(n9775) );
  XOR2X1_RVT U10526 ( .A1(key[90]), .A2(state[90]), .Y(n9877) );
  XOR2X1_RVT U10527 ( .A1(key[91]), .A2(state[91]), .Y(n9811) );
  OR2X1_RVT U10528 ( .A1(n12864), .A2(n12254), .Y(n9751) );
  XOR2X1_RVT U10529 ( .A1(key[93]), .A2(state[93]), .Y(n9737) );
  XOR2X1_RVT U10530 ( .A1(key[94]), .A2(state[94]), .Y(n9773) );
  OR2X1_RVT U10531 ( .A1(n12854), .A2(n12252), .Y(n9977) );
  XOR2X1_RVT U10532 ( .A1(key[88]), .A2(state[88]), .Y(n9752) );
  XOR2X1_RVT U10533 ( .A1(key[89]), .A2(state[89]), .Y(n9862) );
  XOR2X1_RVT U10534 ( .A1(key[95]), .A2(state[95]), .Y(n9746) );
  AND4X1_RVT U10535 ( .A1(n10519), .A2(n10520), .A3(n10521), .A4(n10522), .Y(
        n10518) );
  AND4X1_RVT U10536 ( .A1(n10523), .A2(n10524), .A3(n10525), .A4(n10526), .Y(
        n10522) );
  AND4X1_RVT U10537 ( .A1(n10527), .A2(n10528), .A3(n10529), .A4(n10530), .Y(
        n10526) );
  OR2X1_RVT U10538 ( .A1(n12240), .A2(n10532), .Y(n10525) );
  OR2X1_RVT U10539 ( .A1(n10533), .A2(n10534), .Y(n10523) );
  OR2X1_RVT U10540 ( .A1(n12848), .A2(n10535), .Y(n10534) );
  AND4X1_RVT U10541 ( .A1(n10536), .A2(n10537), .A3(n10538), .A4(n10539), .Y(
        n10521) );
  OR2X1_RVT U10542 ( .A1(n10540), .A2(n12846), .Y(n10539) );
  AND2X1_RVT U10543 ( .A1(n10541), .A2(n10542), .Y(n10540) );
  AND2X1_RVT U10544 ( .A1(n10543), .A2(n10544), .Y(n10538) );
  OR2X1_RVT U10545 ( .A1(n10545), .A2(n116), .Y(n10544) );
  AND2X1_RVT U10546 ( .A1(n10546), .A2(n10547), .Y(n10545) );
  OR2X1_RVT U10547 ( .A1(n12231), .A2(n10549), .Y(n10547) );
  OR2X1_RVT U10548 ( .A1(n10535), .A2(n10550), .Y(n10546) );
  OR2X1_RVT U10549 ( .A1(n10551), .A2(n12237), .Y(n10543) );
  AND2X1_RVT U10550 ( .A1(n10553), .A2(n10554), .Y(n10551) );
  OR2X1_RVT U10551 ( .A1(n10555), .A2(n10556), .Y(n10537) );
  AND2X1_RVT U10552 ( .A1(n10557), .A2(n10558), .Y(n10555) );
  OR2X1_RVT U10553 ( .A1(n12232), .A2(n10559), .Y(n10558) );
  AND2X1_RVT U10554 ( .A1(n10560), .A2(n10561), .Y(n10557) );
  AND2X1_RVT U10555 ( .A1(n10562), .A2(n10563), .Y(n10536) );
  OR2X1_RVT U10556 ( .A1(n10564), .A2(n12214), .Y(n10563) );
  AND2X1_RVT U10557 ( .A1(n10566), .A2(n10567), .Y(n10564) );
  OR2X1_RVT U10558 ( .A1(n10568), .A2(n10569), .Y(n10567) );
  OR2X1_RVT U10559 ( .A1(n12223), .A2(n12218), .Y(n10569) );
  OR2X1_RVT U10560 ( .A1(n10572), .A2(n10573), .Y(n10562) );
  AND2X1_RVT U10561 ( .A1(n10574), .A2(n10575), .Y(n10572) );
  AND2X1_RVT U10562 ( .A1(n10576), .A2(n10577), .Y(n10574) );
  AND4X1_RVT U10563 ( .A1(n10578), .A2(n10579), .A3(n10580), .A4(n10581), .Y(
        n10520) );
  AND4X1_RVT U10564 ( .A1(n10582), .A2(n10583), .A3(n10584), .A4(n10585), .Y(
        n10581) );
  OR2X1_RVT U10565 ( .A1(n10586), .A2(n12243), .Y(n10585) );
  AND4X1_RVT U10566 ( .A1(n10588), .A2(n10589), .A3(n10590), .A4(n10591), .Y(
        n10586) );
  OR2X1_RVT U10567 ( .A1(n10592), .A2(n10559), .Y(n10591) );
  OR2X1_RVT U10568 ( .A1(n10593), .A2(n12229), .Y(n10590) );
  OR2X1_RVT U10569 ( .A1(n10595), .A2(n12220), .Y(n10584) );
  AND4X1_RVT U10570 ( .A1(n10596), .A2(n10597), .A3(n10598), .A4(n10599), .Y(
        n10595) );
  OR2X1_RVT U10571 ( .A1(n10600), .A2(n10601), .Y(n10599) );
  OR2X1_RVT U10572 ( .A1(n12237), .A2(n12232), .Y(n10601) );
  AND2X1_RVT U10573 ( .A1(n10602), .A2(n10603), .Y(n10598) );
  OR2X1_RVT U10574 ( .A1(n12850), .A2(n10604), .Y(n10597) );
  OR2X1_RVT U10575 ( .A1(n10605), .A2(n10606), .Y(n10596) );
  AND2X1_RVT U10576 ( .A1(n10607), .A2(n10608), .Y(n10605) );
  OR2X1_RVT U10577 ( .A1(n12237), .A2(n10609), .Y(n10608) );
  OR2X1_RVT U10578 ( .A1(n10542), .A2(n10610), .Y(n10583) );
  OR2X1_RVT U10579 ( .A1(n10609), .A2(n10611), .Y(n10582) );
  OR2X1_RVT U10580 ( .A1(n10612), .A2(n10613), .Y(n10580) );
  OR2X1_RVT U10581 ( .A1(n10614), .A2(n10607), .Y(n10579) );
  OR2X1_RVT U10582 ( .A1(n10615), .A2(n10616), .Y(n10578) );
  AND4X1_RVT U10583 ( .A1(n10617), .A2(n10618), .A3(n10619), .A4(n10620), .Y(
        n10519) );
  AND2X1_RVT U10584 ( .A1(n10621), .A2(n10622), .Y(n10620) );
  OR2X1_RVT U10585 ( .A1(n10606), .A2(n10623), .Y(n10622) );
  AND2X1_RVT U10586 ( .A1(n10624), .A2(n10625), .Y(n10621) );
  OR2X1_RVT U10587 ( .A1(n10626), .A2(n10549), .Y(n10625) );
  OR2X1_RVT U10588 ( .A1(n10550), .A2(n10627), .Y(n10624) );
  OR2X1_RVT U10589 ( .A1(n114), .A2(n10628), .Y(n10619) );
  OR2X1_RVT U10590 ( .A1(n10629), .A2(n12227), .Y(n10618) );
  OR2X1_RVT U10591 ( .A1(n12230), .A2(n10631), .Y(n10617) );
  AND4X1_RVT U10592 ( .A1(n10633), .A2(n10634), .A3(n10635), .A4(n10636), .Y(
        n10632) );
  AND4X1_RVT U10593 ( .A1(n10637), .A2(n10528), .A3(n10638), .A4(n10639), .Y(
        n10636) );
  AND4X1_RVT U10594 ( .A1(n10640), .A2(n10641), .A3(n10642), .A4(n10643), .Y(
        n10639) );
  OR2X1_RVT U10595 ( .A1(n10549), .A2(n10644), .Y(n10643) );
  OR2X1_RVT U10596 ( .A1(n10645), .A2(n12242), .Y(n10644) );
  OR2X1_RVT U10597 ( .A1(n10550), .A2(n10646), .Y(n10642) );
  OR2X1_RVT U10598 ( .A1(n114), .A2(n12226), .Y(n10646) );
  OR2X1_RVT U10599 ( .A1(n10647), .A2(n10593), .Y(n10641) );
  AND2X1_RVT U10600 ( .A1(n10604), .A2(n10648), .Y(n10647) );
  OR2X1_RVT U10601 ( .A1(n10649), .A2(n10650), .Y(n10640) );
  AND2X1_RVT U10602 ( .A1(n10651), .A2(n10652), .Y(n10649) );
  AND2X1_RVT U10603 ( .A1(n10653), .A2(n10654), .Y(n10638) );
  OR2X1_RVT U10604 ( .A1(n10600), .A2(n10655), .Y(n10654) );
  OR2X1_RVT U10605 ( .A1(n10656), .A2(n12848), .Y(n10655) );
  OR2X1_RVT U10606 ( .A1(n10657), .A2(n10658), .Y(n10653) );
  OR2X1_RVT U10607 ( .A1(n10659), .A2(n12231), .Y(n10658) );
  OR2X1_RVT U10608 ( .A1(n10535), .A2(n10660), .Y(n10528) );
  AND4X1_RVT U10609 ( .A1(n10661), .A2(n10662), .A3(n10663), .A4(n10664), .Y(
        n10635) );
  AND4X1_RVT U10610 ( .A1(n10665), .A2(n10666), .A3(n10667), .A4(n10668), .Y(
        n10664) );
  OR2X1_RVT U10611 ( .A1(n10669), .A2(n12245), .Y(n10668) );
  AND2X1_RVT U10612 ( .A1(n10671), .A2(n10672), .Y(n10669) );
  OR2X1_RVT U10613 ( .A1(n12214), .A2(n10550), .Y(n10672) );
  OR2X1_RVT U10614 ( .A1(n10673), .A2(n10552), .Y(n10667) );
  AND2X1_RVT U10615 ( .A1(n10674), .A2(n10675), .Y(n10673) );
  OR2X1_RVT U10616 ( .A1(n10676), .A2(n12847), .Y(n10666) );
  AND2X1_RVT U10617 ( .A1(n10677), .A2(n10678), .Y(n10676) );
  OR2X1_RVT U10618 ( .A1(n10679), .A2(n10628), .Y(n10678) );
  AND2X1_RVT U10619 ( .A1(n12245), .A2(n12229), .Y(n10679) );
  OR2X1_RVT U10620 ( .A1(n10680), .A2(n12215), .Y(n10665) );
  AND2X1_RVT U10621 ( .A1(n10682), .A2(n10683), .Y(n10680) );
  OR2X1_RVT U10622 ( .A1(n10684), .A2(n12221), .Y(n10663) );
  AND2X1_RVT U10623 ( .A1(n10685), .A2(n10686), .Y(n10684) );
  OR2X1_RVT U10624 ( .A1(n12229), .A2(n10687), .Y(n10686) );
  AND2X1_RVT U10625 ( .A1(n10688), .A2(n10689), .Y(n10685) );
  OR2X1_RVT U10626 ( .A1(n10690), .A2(n10691), .Y(n10688) );
  OR2X1_RVT U10627 ( .A1(n10535), .A2(n10606), .Y(n10691) );
  OR2X1_RVT U10628 ( .A1(n10692), .A2(n12844), .Y(n10662) );
  AND2X1_RVT U10629 ( .A1(n10693), .A2(n10694), .Y(n10692) );
  OR2X1_RVT U10630 ( .A1(n10695), .A2(n10696), .Y(n10661) );
  AND2X1_RVT U10631 ( .A1(n10697), .A2(n10698), .Y(n10695) );
  AND2X1_RVT U10632 ( .A1(n10699), .A2(n10700), .Y(n10697) );
  OR2X1_RVT U10633 ( .A1(n116), .A2(n10628), .Y(n10700) );
  OR2X1_RVT U10634 ( .A1(n12239), .A2(n10593), .Y(n10699) );
  AND4X1_RVT U10635 ( .A1(n10701), .A2(n10702), .A3(n10703), .A4(n10704), .Y(
        n10634) );
  AND4X1_RVT U10636 ( .A1(n10705), .A2(n10706), .A3(n10707), .A4(n10708), .Y(
        n10704) );
  OR2X1_RVT U10637 ( .A1(n10628), .A2(n10627), .Y(n10708) );
  OR2X1_RVT U10638 ( .A1(n10559), .A2(n10709), .Y(n10707) );
  OR2X1_RVT U10639 ( .A1(n10592), .A2(n10710), .Y(n10706) );
  OR2X1_RVT U10640 ( .A1(n10535), .A2(n10711), .Y(n10705) );
  AND2X1_RVT U10641 ( .A1(n10712), .A2(n10713), .Y(n10703) );
  OR2X1_RVT U10642 ( .A1(n12240), .A2(n10714), .Y(n10713) );
  OR2X1_RVT U10643 ( .A1(n12219), .A2(n10611), .Y(n10712) );
  OR2X1_RVT U10644 ( .A1(n10715), .A2(n10570), .Y(n10702) );
  AND4X1_RVT U10645 ( .A1(n10716), .A2(n10717), .A3(n10718), .A4(n10719), .Y(
        n10715) );
  OR2X1_RVT U10646 ( .A1(n10720), .A2(n10535), .Y(n10718) );
  OR2X1_RVT U10647 ( .A1(n12836), .A2(n10721), .Y(n10717) );
  OR2X1_RVT U10648 ( .A1(n10722), .A2(n12844), .Y(n10716) );
  AND2X1_RVT U10649 ( .A1(n10613), .A2(n10723), .Y(n10722) );
  OR2X1_RVT U10650 ( .A1(n10615), .A2(n10724), .Y(n10701) );
  AND4X1_RVT U10651 ( .A1(n10725), .A2(n10726), .A3(n10727), .A4(n10728), .Y(
        n10633) );
  AND4X1_RVT U10652 ( .A1(n10729), .A2(n10730), .A3(n10731), .A4(n10732), .Y(
        n10728) );
  OR2X1_RVT U10653 ( .A1(n12840), .A2(n10733), .Y(n10732) );
  OR2X1_RVT U10654 ( .A1(n12841), .A2(n10734), .Y(n10731) );
  OR2X1_RVT U10655 ( .A1(n12838), .A2(n10735), .Y(n10730) );
  OR2X1_RVT U10656 ( .A1(n12213), .A2(n10736), .Y(n10729) );
  OR2X1_RVT U10657 ( .A1(n10737), .A2(n12220), .Y(n10726) );
  AND4X1_RVT U10658 ( .A1(n10739), .A2(n10740), .A3(n10741), .A4(n10742), .Y(
        n10738) );
  AND4X1_RVT U10659 ( .A1(n10743), .A2(n10744), .A3(n10745), .A4(n10746), .Y(
        n10742) );
  AND4X1_RVT U10660 ( .A1(n10747), .A2(n10524), .A3(n10694), .A4(n10748), .Y(
        n10746) );
  OR2X1_RVT U10661 ( .A1(n10749), .A2(n12835), .Y(n10524) );
  AND2X1_RVT U10662 ( .A1(n10750), .A2(n10751), .Y(n10749) );
  OR2X1_RVT U10663 ( .A1(n10568), .A2(n10752), .Y(n10751) );
  OR2X1_RVT U10664 ( .A1(n10753), .A2(n10650), .Y(n10750) );
  OR2X1_RVT U10665 ( .A1(n10754), .A2(n10609), .Y(n10747) );
  AND2X1_RVT U10666 ( .A1(n10755), .A2(n10756), .Y(n10754) );
  OR2X1_RVT U10667 ( .A1(n12840), .A2(n10593), .Y(n10756) );
  OR2X1_RVT U10668 ( .A1(n10757), .A2(n10552), .Y(n10745) );
  AND2X1_RVT U10669 ( .A1(n10758), .A2(n10759), .Y(n10757) );
  OR2X1_RVT U10670 ( .A1(n10760), .A2(n12846), .Y(n10759) );
  AND2X1_RVT U10671 ( .A1(n10600), .A2(n10761), .Y(n10760) );
  OR2X1_RVT U10672 ( .A1(n10762), .A2(n12240), .Y(n10744) );
  AND2X1_RVT U10673 ( .A1(n10763), .A2(n10764), .Y(n10762) );
  OR2X1_RVT U10674 ( .A1(n10593), .A2(n10559), .Y(n10764) );
  OR2X1_RVT U10675 ( .A1(n10765), .A2(n12223), .Y(n10743) );
  AND2X1_RVT U10676 ( .A1(n10677), .A2(n10766), .Y(n10765) );
  OR2X1_RVT U10677 ( .A1(n10606), .A2(n10767), .Y(n10677) );
  AND4X1_RVT U10678 ( .A1(n10768), .A2(n10769), .A3(n10770), .A4(n10771), .Y(
        n10741) );
  OR2X1_RVT U10679 ( .A1(n10772), .A2(n12230), .Y(n10771) );
  AND2X1_RVT U10680 ( .A1(n10773), .A2(n10774), .Y(n10772) );
  OR2X1_RVT U10681 ( .A1(n10650), .A2(n10550), .Y(n10774) );
  AND2X1_RVT U10682 ( .A1(n10775), .A2(n10776), .Y(n10773) );
  OR2X1_RVT U10683 ( .A1(n10690), .A2(n10752), .Y(n10775) );
  AND2X1_RVT U10684 ( .A1(n10777), .A2(n10778), .Y(n10770) );
  OR2X1_RVT U10685 ( .A1(n10779), .A2(n10681), .Y(n10778) );
  AND2X1_RVT U10686 ( .A1(n10780), .A2(n10589), .Y(n10779) );
  OR2X1_RVT U10687 ( .A1(n10535), .A2(n10650), .Y(n10589) );
  OR2X1_RVT U10688 ( .A1(n10781), .A2(n116), .Y(n10777) );
  AND2X1_RVT U10689 ( .A1(n10782), .A2(n10783), .Y(n10781) );
  OR2X1_RVT U10690 ( .A1(n10784), .A2(n12232), .Y(n10783) );
  AND2X1_RVT U10691 ( .A1(n10785), .A2(n10786), .Y(n10784) );
  OR2X1_RVT U10692 ( .A1(n12227), .A2(n10600), .Y(n10786) );
  OR2X1_RVT U10693 ( .A1(n12850), .A2(n12229), .Y(n10785) );
  AND2X1_RVT U10694 ( .A1(n10651), .A2(n10761), .Y(n10782) );
  OR2X1_RVT U10695 ( .A1(n10681), .A2(n10787), .Y(n10651) );
  OR2X1_RVT U10696 ( .A1(n12845), .A2(n12841), .Y(n10787) );
  OR2X1_RVT U10697 ( .A1(n10788), .A2(n10670), .Y(n10769) );
  AND4X1_RVT U10698 ( .A1(n10629), .A2(n10789), .A3(n10790), .A4(n10791), .Y(
        n10788) );
  OR2X1_RVT U10699 ( .A1(n12231), .A2(n10650), .Y(n10791) );
  AND2X1_RVT U10700 ( .A1(n10792), .A2(n10793), .Y(n10790) );
  OR2X1_RVT U10701 ( .A1(n12850), .A2(n12240), .Y(n10789) );
  AND2X1_RVT U10702 ( .A1(n10794), .A2(n10795), .Y(n10629) );
  OR2X1_RVT U10703 ( .A1(n10796), .A2(n114), .Y(n10795) );
  OR2X1_RVT U10704 ( .A1(n10593), .A2(n12835), .Y(n10794) );
  AND2X1_RVT U10705 ( .A1(n10797), .A2(n10798), .Y(n10768) );
  OR2X1_RVT U10706 ( .A1(n10799), .A2(n12837), .Y(n10798) );
  AND2X1_RVT U10707 ( .A1(n10800), .A2(n10801), .Y(n10799) );
  OR2X1_RVT U10708 ( .A1(n10802), .A2(n12234), .Y(n10801) );
  AND2X1_RVT U10709 ( .A1(n10803), .A2(n10804), .Y(n10802) );
  AND2X1_RVT U10710 ( .A1(n10805), .A2(n10806), .Y(n10800) );
  OR2X1_RVT U10711 ( .A1(n10807), .A2(n12243), .Y(n10797) );
  AND4X1_RVT U10712 ( .A1(n10808), .A2(n10809), .A3(n10810), .A4(n10811), .Y(
        n10807) );
  OR2X1_RVT U10713 ( .A1(n12849), .A2(n10812), .Y(n10810) );
  OR2X1_RVT U10714 ( .A1(n114), .A2(n10607), .Y(n10809) );
  OR2X1_RVT U10715 ( .A1(n10696), .A2(n10650), .Y(n10808) );
  AND4X1_RVT U10716 ( .A1(n10813), .A2(n10814), .A3(n10815), .A4(n10816), .Y(
        n10740) );
  AND2X1_RVT U10717 ( .A1(n10817), .A2(n10660), .Y(n10816) );
  OR2X1_RVT U10718 ( .A1(n12218), .A2(n10626), .Y(n10660) );
  AND2X1_RVT U10719 ( .A1(n10818), .A2(n10819), .Y(n10817) );
  OR2X1_RVT U10720 ( .A1(n10820), .A2(n10575), .Y(n10819) );
  OR2X1_RVT U10721 ( .A1(n10627), .A2(n10687), .Y(n10818) );
  OR2X1_RVT U10722 ( .A1(n114), .A2(n10821), .Y(n10815) );
  OR2X1_RVT U10723 ( .A1(n12848), .A2(n10822), .Y(n10814) );
  OR2X1_RVT U10724 ( .A1(n10696), .A2(n10823), .Y(n10813) );
  AND4X1_RVT U10725 ( .A1(n10824), .A2(n10825), .A3(n10826), .A4(n10827), .Y(
        n10739) );
  AND2X1_RVT U10726 ( .A1(n10828), .A2(n10829), .Y(n10827) );
  OR2X1_RVT U10727 ( .A1(n12213), .A2(n10830), .Y(n10829) );
  AND2X1_RVT U10728 ( .A1(n10831), .A2(n10832), .Y(n10828) );
  OR2X1_RVT U10729 ( .A1(n10592), .A2(n10602), .Y(n10832) );
  OR2X1_RVT U10730 ( .A1(n12234), .A2(n10652), .Y(n10602) );
  OR2X1_RVT U10731 ( .A1(n12220), .A2(n10833), .Y(n10831) );
  OR2X1_RVT U10732 ( .A1(n10573), .A2(n10566), .Y(n10826) );
  OR2X1_RVT U10733 ( .A1(n10659), .A2(n10834), .Y(n10566) );
  OR2X1_RVT U10734 ( .A1(n12844), .A2(n10835), .Y(n10825) );
  OR2X1_RVT U10735 ( .A1(n12232), .A2(n10693), .Y(n10824) );
  OR2X1_RVT U10736 ( .A1(n12835), .A2(n10755), .Y(n10693) );
  AND4X1_RVT U10737 ( .A1(n10837), .A2(n10838), .A3(n10839), .A4(n10840), .Y(
        n10836) );
  AND4X1_RVT U10738 ( .A1(n10841), .A2(n10842), .A3(n10843), .A4(n10844), .Y(
        n10840) );
  OR2X1_RVT U10739 ( .A1(n124), .A2(n10845), .Y(n10844) );
  OR2X1_RVT U10740 ( .A1(n10846), .A2(n12245), .Y(n10845) );
  AND2X1_RVT U10741 ( .A1(n12234), .A2(n10612), .Y(n10846) );
  AND2X1_RVT U10742 ( .A1(n10527), .A2(n10847), .Y(n10843) );
  OR2X1_RVT U10743 ( .A1(n12223), .A2(n10848), .Y(n10527) );
  OR2X1_RVT U10744 ( .A1(n124), .A2(n10606), .Y(n10848) );
  OR2X1_RVT U10745 ( .A1(n10849), .A2(n10535), .Y(n10842) );
  AND2X1_RVT U10746 ( .A1(n10850), .A2(n10851), .Y(n10849) );
  AND2X1_RVT U10747 ( .A1(n10852), .A2(n10853), .Y(n10841) );
  OR2X1_RVT U10748 ( .A1(n10854), .A2(n10855), .Y(n10853) );
  AND2X1_RVT U10749 ( .A1(n10856), .A2(n10616), .Y(n10854) );
  OR2X1_RVT U10750 ( .A1(n10857), .A2(n10607), .Y(n10852) );
  AND2X1_RVT U10751 ( .A1(n10792), .A2(n10626), .Y(n10857) );
  OR2X1_RVT U10752 ( .A1(n12221), .A2(n10858), .Y(n10792) );
  OR2X1_RVT U10753 ( .A1(n12850), .A2(n12231), .Y(n10858) );
  AND4X1_RVT U10754 ( .A1(n10859), .A2(n10860), .A3(n10861), .A4(n10862), .Y(
        n10839) );
  OR2X1_RVT U10755 ( .A1(n10863), .A2(n12840), .Y(n10862) );
  AND2X1_RVT U10756 ( .A1(n10675), .A2(n10864), .Y(n10863) );
  OR2X1_RVT U10757 ( .A1(n12848), .A2(n10720), .Y(n10675) );
  AND2X1_RVT U10758 ( .A1(n10865), .A2(n10866), .Y(n10861) );
  OR2X1_RVT U10759 ( .A1(n10867), .A2(n12838), .Y(n10866) );
  AND2X1_RVT U10760 ( .A1(n10868), .A2(n10869), .Y(n10867) );
  OR2X1_RVT U10761 ( .A1(n10570), .A2(n10812), .Y(n10869) );
  OR2X1_RVT U10762 ( .A1(n10870), .A2(n12836), .Y(n10865) );
  AND2X1_RVT U10763 ( .A1(n10871), .A2(n10872), .Y(n10870) );
  OR2X1_RVT U10764 ( .A1(n10873), .A2(n12234), .Y(n10860) );
  AND2X1_RVT U10765 ( .A1(n10874), .A2(n10875), .Y(n10873) );
  AND2X1_RVT U10766 ( .A1(n10876), .A2(n10877), .Y(n10874) );
  AND2X1_RVT U10767 ( .A1(n10878), .A2(n10879), .Y(n10859) );
  OR2X1_RVT U10768 ( .A1(n10880), .A2(n10796), .Y(n10879) );
  AND2X1_RVT U10769 ( .A1(n10881), .A2(n10627), .Y(n10880) );
  AND2X1_RVT U10770 ( .A1(n10882), .A2(n10883), .Y(n10881) );
  OR2X1_RVT U10771 ( .A1(n10884), .A2(n12237), .Y(n10878) );
  AND2X1_RVT U10772 ( .A1(n10885), .A2(n10886), .Y(n10884) );
  OR2X1_RVT U10773 ( .A1(n12847), .A2(n12239), .Y(n10886) );
  AND2X1_RVT U10774 ( .A1(n10616), .A2(n10887), .Y(n10885) );
  AND4X1_RVT U10775 ( .A1(n10888), .A2(n10889), .A3(n10890), .A4(n10891), .Y(
        n10838) );
  AND2X1_RVT U10776 ( .A1(n10892), .A2(n10893), .Y(n10891) );
  OR2X1_RVT U10777 ( .A1(n10609), .A2(n10683), .Y(n10893) );
  OR2X1_RVT U10778 ( .A1(n12842), .A2(n10616), .Y(n10683) );
  AND2X1_RVT U10779 ( .A1(n10894), .A2(n10895), .Y(n10892) );
  OR2X1_RVT U10780 ( .A1(n10761), .A2(n10575), .Y(n10895) );
  OR2X1_RVT U10781 ( .A1(n12849), .A2(n12230), .Y(n10575) );
  OR2X1_RVT U10782 ( .A1(n10659), .A2(n10709), .Y(n10894) );
  OR2X1_RVT U10783 ( .A1(n12837), .A2(n10896), .Y(n10709) );
  OR2X1_RVT U10784 ( .A1(n10897), .A2(n12213), .Y(n10890) );
  AND4X1_RVT U10785 ( .A1(n10898), .A2(n10899), .A3(n10900), .A4(n10901), .Y(
        n10897) );
  OR2X1_RVT U10786 ( .A1(n10834), .A2(n10607), .Y(n10900) );
  OR2X1_RVT U10787 ( .A1(n10902), .A2(n10604), .Y(n10899) );
  OR2X1_RVT U10788 ( .A1(n12846), .A2(n10559), .Y(n10898) );
  OR2X1_RVT U10789 ( .A1(n10903), .A2(n12214), .Y(n10889) );
  AND2X1_RVT U10790 ( .A1(n10904), .A2(n10905), .Y(n10903) );
  OR2X1_RVT U10791 ( .A1(n10834), .A2(n10559), .Y(n10905) );
  AND2X1_RVT U10792 ( .A1(n10906), .A2(n10835), .Y(n10904) );
  OR2X1_RVT U10793 ( .A1(n10607), .A2(n10907), .Y(n10835) );
  OR2X1_RVT U10794 ( .A1(n12837), .A2(n12849), .Y(n10907) );
  OR2X1_RVT U10795 ( .A1(n10908), .A2(n12221), .Y(n10888) );
  AND4X1_RVT U10796 ( .A1(n10909), .A2(n10822), .A3(n10631), .A4(n10603), .Y(
        n10908) );
  OR2X1_RVT U10797 ( .A1(n10628), .A2(n10910), .Y(n10603) );
  OR2X1_RVT U10798 ( .A1(n12839), .A2(n10565), .Y(n10910) );
  OR2X1_RVT U10799 ( .A1(n10690), .A2(n10724), .Y(n10631) );
  OR2X1_RVT U10800 ( .A1(n10609), .A2(n10911), .Y(n10822) );
  OR2X1_RVT U10801 ( .A1(n12245), .A2(n12214), .Y(n10911) );
  OR2X1_RVT U10802 ( .A1(n10568), .A2(n10912), .Y(n10909) );
  OR2X1_RVT U10803 ( .A1(n10913), .A2(n12219), .Y(n10912) );
  AND4X1_RVT U10804 ( .A1(n10914), .A2(n10915), .A3(n10916), .A4(n10917), .Y(
        n10837) );
  AND2X1_RVT U10805 ( .A1(n10918), .A2(n10919), .Y(n10917) );
  AND2X1_RVT U10806 ( .A1(n10920), .A2(n10921), .Y(n10918) );
  OR2X1_RVT U10807 ( .A1(n10600), .A2(n10875), .Y(n10921) );
  OR2X1_RVT U10808 ( .A1(n10612), .A2(n10922), .Y(n10875) );
  OR2X1_RVT U10809 ( .A1(n12838), .A2(n12840), .Y(n10922) );
  OR2X1_RVT U10810 ( .A1(n12845), .A2(n10923), .Y(n10920) );
  OR2X1_RVT U10811 ( .A1(n12230), .A2(n10924), .Y(n10916) );
  OR2X1_RVT U10812 ( .A1(n12848), .A2(n10925), .Y(n10915) );
  OR2X1_RVT U10813 ( .A1(n10612), .A2(n10926), .Y(n10914) );
  AND4X1_RVT U10814 ( .A1(n10928), .A2(n10929), .A3(n10930), .A4(n10931), .Y(
        n10927) );
  AND4X1_RVT U10815 ( .A1(n10932), .A2(n10933), .A3(n10934), .A4(n10935), .Y(
        n10931) );
  AND4X1_RVT U10816 ( .A1(n10936), .A2(n10937), .A3(n10529), .A4(n10938), .Y(
        n10935) );
  OR2X1_RVT U10817 ( .A1(n10670), .A2(n10939), .Y(n10529) );
  OR2X1_RVT U10818 ( .A1(n10761), .A2(n116), .Y(n10939) );
  OR2X1_RVT U10819 ( .A1(n10533), .A2(n10940), .Y(n10937) );
  OR2X1_RVT U10820 ( .A1(n12843), .A2(n12846), .Y(n10940) );
  OR2X1_RVT U10821 ( .A1(n10796), .A2(n10941), .Y(n10936) );
  OR2X1_RVT U10822 ( .A1(n10942), .A2(n10570), .Y(n10941) );
  AND2X1_RVT U10823 ( .A1(n12234), .A2(n10670), .Y(n10942) );
  OR2X1_RVT U10824 ( .A1(n10943), .A2(n12240), .Y(n10934) );
  AND2X1_RVT U10825 ( .A1(n10811), .A2(n10883), .Y(n10943) );
  OR2X1_RVT U10826 ( .A1(n116), .A2(n10944), .Y(n10883) );
  OR2X1_RVT U10827 ( .A1(n12213), .A2(n12842), .Y(n10944) );
  OR2X1_RVT U10828 ( .A1(n10600), .A2(n10945), .Y(n10811) );
  OR2X1_RVT U10829 ( .A1(n12840), .A2(n10592), .Y(n10945) );
  OR2X1_RVT U10830 ( .A1(n10946), .A2(n10550), .Y(n10933) );
  AND2X1_RVT U10831 ( .A1(n10947), .A2(n10755), .Y(n10946) );
  OR2X1_RVT U10832 ( .A1(n10656), .A2(n10650), .Y(n10932) );
  AND4X1_RVT U10833 ( .A1(n10948), .A2(n10949), .A3(n10950), .A4(n10951), .Y(
        n10930) );
  AND2X1_RVT U10834 ( .A1(n10952), .A2(n10953), .Y(n10951) );
  OR2X1_RVT U10835 ( .A1(n10954), .A2(n12234), .Y(n10953) );
  AND2X1_RVT U10836 ( .A1(n10955), .A2(n10623), .Y(n10954) );
  AND2X1_RVT U10837 ( .A1(n10956), .A2(n10957), .Y(n10952) );
  OR2X1_RVT U10838 ( .A1(n10958), .A2(n10606), .Y(n10957) );
  AND2X1_RVT U10839 ( .A1(n10577), .A2(n10549), .Y(n10958) );
  OR2X1_RVT U10840 ( .A1(n12848), .A2(n10648), .Y(n10577) );
  OR2X1_RVT U10841 ( .A1(n10959), .A2(n10659), .Y(n10956) );
  AND2X1_RVT U10842 ( .A1(n10851), .A2(n10960), .Y(n10959) );
  OR2X1_RVT U10843 ( .A1(n12849), .A2(n10687), .Y(n10851) );
  OR2X1_RVT U10844 ( .A1(n10961), .A2(n12840), .Y(n10950) );
  AND2X1_RVT U10845 ( .A1(n10554), .A2(n10962), .Y(n10961) );
  OR2X1_RVT U10846 ( .A1(n10690), .A2(n10614), .Y(n10962) );
  OR2X1_RVT U10847 ( .A1(n10593), .A2(n10796), .Y(n10554) );
  OR2X1_RVT U10848 ( .A1(n10963), .A2(n114), .Y(n10949) );
  AND2X1_RVT U10849 ( .A1(n10604), .A2(n10964), .Y(n10963) );
  OR2X1_RVT U10850 ( .A1(n10965), .A2(n12218), .Y(n10964) );
  AND2X1_RVT U10851 ( .A1(n10966), .A2(n10967), .Y(n10965) );
  OR2X1_RVT U10852 ( .A1(n12841), .A2(n10587), .Y(n10967) );
  OR2X1_RVT U10853 ( .A1(n12245), .A2(n10690), .Y(n10604) );
  OR2X1_RVT U10854 ( .A1(n10968), .A2(n10674), .Y(n10948) );
  AND2X1_RVT U10855 ( .A1(n10607), .A2(n10652), .Y(n10968) );
  OR2X1_RVT U10856 ( .A1(n12837), .A2(n10535), .Y(n10652) );
  AND4X1_RVT U10857 ( .A1(n10969), .A2(n10970), .A3(n10971), .A4(n10972), .Y(
        n10929) );
  AND4X1_RVT U10858 ( .A1(n10973), .A2(n10974), .A3(n10975), .A4(n10976), .Y(
        n10972) );
  OR2X1_RVT U10859 ( .A1(n10977), .A2(n12848), .Y(n10976) );
  AND2X1_RVT U10860 ( .A1(n10710), .A2(n10978), .Y(n10977) );
  OR2X1_RVT U10861 ( .A1(n12242), .A2(n10559), .Y(n10978) );
  OR2X1_RVT U10862 ( .A1(n10979), .A2(n10552), .Y(n10975) );
  AND2X1_RVT U10863 ( .A1(n10980), .A2(n10981), .Y(n10979) );
  OR2X1_RVT U10864 ( .A1(n10982), .A2(n10587), .Y(n10981) );
  AND2X1_RVT U10865 ( .A1(n10612), .A2(n10600), .Y(n10982) );
  AND2X1_RVT U10866 ( .A1(n10614), .A2(n10856), .Y(n10980) );
  OR2X1_RVT U10867 ( .A1(n12243), .A2(n10752), .Y(n10856) );
  OR2X1_RVT U10868 ( .A1(n10983), .A2(n12232), .Y(n10974) );
  AND2X1_RVT U10869 ( .A1(n10984), .A2(n10985), .Y(n10983) );
  OR2X1_RVT U10870 ( .A1(n10600), .A2(n10986), .Y(n10985) );
  AND2X1_RVT U10871 ( .A1(n10682), .A2(n10876), .Y(n10984) );
  OR2X1_RVT U10872 ( .A1(n10592), .A2(n10767), .Y(n10876) );
  OR2X1_RVT U10873 ( .A1(n10565), .A2(n10987), .Y(n10682) );
  OR2X1_RVT U10874 ( .A1(n10988), .A2(n10535), .Y(n10973) );
  AND4X1_RVT U10875 ( .A1(n10989), .A2(n10990), .A3(n10991), .A4(n10924), .Y(
        n10988) );
  OR2X1_RVT U10876 ( .A1(n10628), .A2(n10992), .Y(n10924) );
  OR2X1_RVT U10877 ( .A1(n12213), .A2(n10592), .Y(n10992) );
  OR2X1_RVT U10878 ( .A1(n12845), .A2(n10834), .Y(n10990) );
  OR2X1_RVT U10879 ( .A1(n10593), .A2(n10690), .Y(n10989) );
  OR2X1_RVT U10880 ( .A1(n10761), .A2(n10803), .Y(n10971) );
  OR2X1_RVT U10881 ( .A1(n10993), .A2(n12216), .Y(n10970) );
  AND4X1_RVT U10882 ( .A1(n10994), .A2(n10995), .A3(n10637), .A4(n10735), .Y(
        n10993) );
  OR2X1_RVT U10883 ( .A1(n10559), .A2(n10724), .Y(n10735) );
  OR2X1_RVT U10884 ( .A1(n12845), .A2(n114), .Y(n10724) );
  OR2X1_RVT U10885 ( .A1(n10552), .A2(n10616), .Y(n10637) );
  OR2X1_RVT U10886 ( .A1(n12837), .A2(n10987), .Y(n10969) );
  AND4X1_RVT U10887 ( .A1(n10996), .A2(n10997), .A3(n10998), .A4(n10999), .Y(
        n10928) );
  OR2X1_RVT U10888 ( .A1(n12221), .A2(n11000), .Y(n10999) );
  AND2X1_RVT U10889 ( .A1(n11001), .A2(n11002), .Y(n10998) );
  OR2X1_RVT U10890 ( .A1(n12242), .A2(n10755), .Y(n11002) );
  OR2X1_RVT U10891 ( .A1(n10542), .A2(n10616), .Y(n11001) );
  OR2X1_RVT U10892 ( .A1(n116), .A2(n10573), .Y(n10616) );
  OR2X1_RVT U10893 ( .A1(n12245), .A2(n10734), .Y(n10997) );
  OR2X1_RVT U10894 ( .A1(n10609), .A2(n11003), .Y(n10734) );
  AND2X1_RVT U10895 ( .A1(n11004), .A2(n11005), .Y(n10996) );
  OR2X1_RVT U10896 ( .A1(n12214), .A2(n11006), .Y(n11005) );
  OR2X1_RVT U10897 ( .A1(n10612), .A2(n10561), .Y(n11004) );
  OR2X1_RVT U10898 ( .A1(n10535), .A2(n10820), .Y(n10561) );
  AND4X1_RVT U10899 ( .A1(n11008), .A2(n11009), .A3(n11010), .A4(n11011), .Y(
        n11007) );
  AND4X1_RVT U10900 ( .A1(n11012), .A2(n11013), .A3(n11014), .A4(n11015), .Y(
        n11011) );
  AND4X1_RVT U10901 ( .A1(n8054), .A2(n10028), .A3(n11016), .A4(n11017), .Y(
        n11015) );
  OR2X1_RVT U10902 ( .A1(n10042), .A2(n6196), .Y(n10028) );
  OR2X1_RVT U10903 ( .A1(n6199), .A2(n11018), .Y(n8054) );
  AND4X1_RVT U10904 ( .A1(n11019), .A2(n8130), .A3(n6965), .A4(n6126), .Y(
        n11014) );
  OR2X1_RVT U10905 ( .A1(n6128), .A2(n11020), .Y(n6126) );
  OR2X1_RVT U10906 ( .A1(n12876), .A2(n12203), .Y(n11020) );
  OR2X1_RVT U10907 ( .A1(n1314), .A2(n11021), .Y(n6965) );
  OR2X1_RVT U10908 ( .A1(n12203), .A2(n1306), .Y(n11021) );
  OR2X1_RVT U10909 ( .A1(n12208), .A2(n11022), .Y(n8130) );
  OR2X1_RVT U10910 ( .A1(n69), .A2(n12189), .Y(n11022) );
  OR2X1_RVT U10911 ( .A1(n1376), .A2(n11023), .Y(n11019) );
  OR2X1_RVT U10912 ( .A1(n8919), .A2(n78), .Y(n11023) );
  OR2X1_RVT U10913 ( .A1(n85), .A2(n12204), .Y(n1376) );
  AND4X1_RVT U10914 ( .A1(n11024), .A2(n11025), .A3(n11026), .A4(n11027), .Y(
        n11013) );
  OR2X1_RVT U10915 ( .A1(n6180), .A2(n8932), .Y(n11027) );
  OR2X1_RVT U10916 ( .A1(n7034), .A2(n1334), .Y(n8932) );
  OR2X1_RVT U10917 ( .A1(n7008), .A2(n11028), .Y(n11026) );
  OR2X1_RVT U10918 ( .A1(n6999), .A2(n8063), .Y(n11028) );
  OR2X1_RVT U10919 ( .A1(n11029), .A2(n6198), .Y(n11025) );
  AND2X1_RVT U10920 ( .A1(n7006), .A2(n11030), .Y(n11029) );
  OR2X1_RVT U10921 ( .A1(n11031), .A2(n12201), .Y(n11024) );
  AND2X1_RVT U10922 ( .A1(n8080), .A2(n8947), .Y(n11031) );
  OR2X1_RVT U10923 ( .A1(n12184), .A2(n1329), .Y(n8947) );
  OR2X1_RVT U10924 ( .A1(n73), .A2(n12869), .Y(n1329) );
  OR2X1_RVT U10925 ( .A1(n73), .A2(n6176), .Y(n8080) );
  OR2X1_RVT U10926 ( .A1(n85), .A2(n12209), .Y(n6176) );
  AND4X1_RVT U10927 ( .A1(n11032), .A2(n11033), .A3(n11034), .A4(n11035), .Y(
        n11012) );
  OR2X1_RVT U10928 ( .A1(n11036), .A2(n1388), .Y(n11035) );
  AND2X1_RVT U10929 ( .A1(n7013), .A2(n11037), .Y(n11036) );
  OR2X1_RVT U10930 ( .A1(n8065), .A2(n11038), .Y(n11037) );
  AND2X1_RVT U10931 ( .A1(n11039), .A2(n11040), .Y(n11038) );
  OR2X1_RVT U10932 ( .A1(n1325), .A2(n12198), .Y(n11039) );
  OR2X1_RVT U10933 ( .A1(n12199), .A2(n12208), .Y(n7013) );
  OR2X1_RVT U10934 ( .A1(n11041), .A2(n12877), .Y(n11034) );
  OR2X1_RVT U10935 ( .A1(n11042), .A2(n85), .Y(n11033) );
  AND2X1_RVT U10936 ( .A1(n11043), .A2(n11044), .Y(n11042) );
  OR2X1_RVT U10937 ( .A1(n8065), .A2(n6199), .Y(n11044) );
  OR2X1_RVT U10938 ( .A1(n12877), .A2(n12201), .Y(n6199) );
  OR2X1_RVT U10939 ( .A1(n76), .A2(n8925), .Y(n11043) );
  OR2X1_RVT U10940 ( .A1(n11045), .A2(n12868), .Y(n11032) );
  AND2X1_RVT U10941 ( .A1(n6156), .A2(n6986), .Y(n11045) );
  OR2X1_RVT U10942 ( .A1(n1314), .A2(n1386), .Y(n6986) );
  OR2X1_RVT U10943 ( .A1(n12872), .A2(n8919), .Y(n1386) );
  OR2X1_RVT U10944 ( .A1(n1314), .A2(n11046), .Y(n6156) );
  OR2X1_RVT U10945 ( .A1(n72), .A2(n12203), .Y(n11046) );
  AND4X1_RVT U10946 ( .A1(n11047), .A2(n11048), .A3(n11049), .A4(n11050), .Y(
        n11010) );
  AND4X1_RVT U10947 ( .A1(n11051), .A2(n11052), .A3(n11053), .A4(n11054), .Y(
        n11050) );
  OR2X1_RVT U10948 ( .A1(n1345), .A2(n8101), .Y(n11054) );
  AND2X1_RVT U10949 ( .A1(n11055), .A2(n1391), .Y(n1345) );
  OR2X1_RVT U10950 ( .A1(n76), .A2(n85), .Y(n11055) );
  OR2X1_RVT U10951 ( .A1(n6200), .A2(n1347), .Y(n11053) );
  OR2X1_RVT U10952 ( .A1(n6132), .A2(n12196), .Y(n1347) );
  OR2X1_RVT U10953 ( .A1(n12192), .A2(n6989), .Y(n11052) );
  OR2X1_RVT U10954 ( .A1(n12198), .A2(n6150), .Y(n11051) );
  OR2X1_RVT U10955 ( .A1(n1314), .A2(n7006), .Y(n6150) );
  OR2X1_RVT U10956 ( .A1(n70), .A2(n12869), .Y(n11049) );
  OR2X1_RVT U10957 ( .A1(n11057), .A2(n11058), .Y(n11056) );
  AND2X1_RVT U10958 ( .A1(n1328), .A2(n8901), .Y(n11058) );
  AND2X1_RVT U10959 ( .A1(n11059), .A2(n8065), .Y(n11057) );
  AND2X1_RVT U10960 ( .A1(n71), .A2(n12874), .Y(n11059) );
  OR2X1_RVT U10961 ( .A1(n72), .A2(n7031), .Y(n11048) );
  OR2X1_RVT U10962 ( .A1(n12185), .A2(n11060), .Y(n7031) );
  OR2X1_RVT U10963 ( .A1(n12211), .A2(n12870), .Y(n11060) );
  OR2X1_RVT U10964 ( .A1(n1300), .A2(n7043), .Y(n11047) );
  OR2X1_RVT U10965 ( .A1(n1332), .A2(n11061), .Y(n7043) );
  OR2X1_RVT U10966 ( .A1(n12926), .A2(n12194), .Y(n11061) );
  AND4X1_RVT U10967 ( .A1(n11062), .A2(n11063), .A3(n11064), .A4(n11065), .Y(
        n11009) );
  OR2X1_RVT U10968 ( .A1(n11066), .A2(n83), .Y(n11065) );
  AND2X1_RVT U10969 ( .A1(n11067), .A2(n11068), .Y(n11066) );
  OR2X1_RVT U10970 ( .A1(n69), .A2(n12195), .Y(n11068) );
  AND2X1_RVT U10971 ( .A1(n11069), .A2(n11070), .Y(n11067) );
  OR2X1_RVT U10972 ( .A1(n12209), .A2(n8101), .Y(n11069) );
  OR2X1_RVT U10973 ( .A1(n12871), .A2(n72), .Y(n8101) );
  OR2X1_RVT U10974 ( .A1(n11071), .A2(n1325), .Y(n11064) );
  AND2X1_RVT U10975 ( .A1(n11072), .A2(n11073), .Y(n11071) );
  OR2X1_RVT U10976 ( .A1(n1306), .A2(n78), .Y(n11073) );
  OR2X1_RVT U10977 ( .A1(n12867), .A2(n12876), .Y(n1306) );
  AND2X1_RVT U10978 ( .A1(n11074), .A2(n8134), .Y(n11072) );
  OR2X1_RVT U10979 ( .A1(n1391), .A2(n6172), .Y(n8134) );
  OR2X1_RVT U10980 ( .A1(n11075), .A2(n6132), .Y(n11063) );
  AND2X1_RVT U10981 ( .A1(n11076), .A2(n6989), .Y(n11075) );
  AND2X1_RVT U10982 ( .A1(n11070), .A2(n7005), .Y(n11076) );
  OR2X1_RVT U10983 ( .A1(n12195), .A2(n8061), .Y(n7005) );
  OR2X1_RVT U10984 ( .A1(n12150), .A2(n11030), .Y(n11070) );
  OR2X1_RVT U10985 ( .A1(n11077), .A2(n12871), .Y(n11062) );
  AND2X1_RVT U10986 ( .A1(n11078), .A2(n10055), .Y(n11077) );
  OR2X1_RVT U10987 ( .A1(n76), .A2(n6180), .Y(n10055) );
  OR2X1_RVT U10988 ( .A1(n12874), .A2(n12870), .Y(n6180) );
  AND2X1_RVT U10989 ( .A1(n7014), .A2(n7049), .Y(n11078) );
  OR2X1_RVT U10990 ( .A1(n1334), .A2(n11079), .Y(n7014) );
  OR2X1_RVT U10991 ( .A1(n69), .A2(n8063), .Y(n11079) );
  AND4X1_RVT U10992 ( .A1(n11080), .A2(n11081), .A3(n11082), .A4(n11083), .Y(
        n11008) );
  OR2X1_RVT U10993 ( .A1(n11084), .A2(n12149), .Y(n11083) );
  AND2X1_RVT U10994 ( .A1(n11085), .A2(n8102), .Y(n11084) );
  OR2X1_RVT U10995 ( .A1(n12870), .A2(n6190), .Y(n8102) );
  OR2X1_RVT U10996 ( .A1(n71), .A2(n1388), .Y(n6190) );
  OR2X1_RVT U10997 ( .A1(n11086), .A2(n8919), .Y(n11085) );
  AND2X1_RVT U10998 ( .A1(n11040), .A2(n11087), .Y(n11086) );
  OR2X1_RVT U10999 ( .A1(n12189), .A2(n1391), .Y(n11087) );
  OR2X1_RVT U11000 ( .A1(n71), .A2(n1332), .Y(n11040) );
  OR2X1_RVT U11001 ( .A1(n6143), .A2(n6196), .Y(n11082) );
  OR2X1_RVT U11002 ( .A1(n8056), .A2(n10073), .Y(n11081) );
  OR2X1_RVT U11003 ( .A1(n12184), .A2(n12192), .Y(n10073) );
  OR2X1_RVT U11004 ( .A1(n7052), .A2(n1390), .Y(n11080) );
  OR2X1_RVT U11005 ( .A1(n12874), .A2(n1300), .Y(n1390) );
  OR2X1_RVT U11006 ( .A1(n12191), .A2(n12209), .Y(n7052) );
  AND4X1_RVT U11007 ( .A1(n11089), .A2(n11090), .A3(n11091), .A4(n11092), .Y(
        n11088) );
  AND4X1_RVT U11008 ( .A1(n11093), .A2(n11094), .A3(n11095), .A4(n11096), .Y(
        n11092) );
  AND4X1_RVT U11009 ( .A1(n10748), .A2(n10938), .A3(n11097), .A4(n11098), .Y(
        n11096) );
  OR2X1_RVT U11010 ( .A1(n11099), .A2(n11100), .Y(n10938) );
  OR2X1_RVT U11011 ( .A1(n10533), .A2(n10803), .Y(n10748) );
  OR2X1_RVT U11012 ( .A1(n12846), .A2(n12230), .Y(n10803) );
  AND4X1_RVT U11013 ( .A1(n11006), .A2(n10872), .A3(n10995), .A4(n10530), .Y(
        n11095) );
  OR2X1_RVT U11014 ( .A1(n11101), .A2(n10720), .Y(n10530) );
  OR2X1_RVT U11015 ( .A1(n10535), .A2(n11102), .Y(n10995) );
  OR2X1_RVT U11016 ( .A1(n10568), .A2(n114), .Y(n10872) );
  OR2X1_RVT U11017 ( .A1(n10559), .A2(n11103), .Y(n11006) );
  OR2X1_RVT U11018 ( .A1(n12220), .A2(n12240), .Y(n11103) );
  AND4X1_RVT U11019 ( .A1(n11104), .A2(n11105), .A3(n11106), .A4(n11107), .Y(
        n11094) );
  OR2X1_RVT U11020 ( .A1(n10812), .A2(n11108), .Y(n11107) );
  OR2X1_RVT U11021 ( .A1(n12240), .A2(n10592), .Y(n11108) );
  OR2X1_RVT U11022 ( .A1(n10721), .A2(n11109), .Y(n11106) );
  OR2X1_RVT U11023 ( .A1(n12847), .A2(n10609), .Y(n11109) );
  OR2X1_RVT U11024 ( .A1(n10947), .A2(n11110), .Y(n11105) );
  OR2X1_RVT U11025 ( .A1(n11111), .A2(n10606), .Y(n11110) );
  OR2X1_RVT U11026 ( .A1(n12237), .A2(n11112), .Y(n11104) );
  OR2X1_RVT U11027 ( .A1(n11113), .A2(n12220), .Y(n11112) );
  AND2X1_RVT U11028 ( .A1(n10820), .A2(n11114), .Y(n11113) );
  AND2X1_RVT U11029 ( .A1(n11115), .A2(n11116), .Y(n11093) );
  OR2X1_RVT U11030 ( .A1(n11117), .A2(n10587), .Y(n11116) );
  AND2X1_RVT U11031 ( .A1(n11118), .A2(n11119), .Y(n11117) );
  OR2X1_RVT U11032 ( .A1(n12219), .A2(n10780), .Y(n11119) );
  OR2X1_RVT U11033 ( .A1(n12223), .A2(n10855), .Y(n11118) );
  AND2X1_RVT U11034 ( .A1(n11120), .A2(n11121), .Y(n11115) );
  OR2X1_RVT U11035 ( .A1(n11122), .A2(n10626), .Y(n11121) );
  AND2X1_RVT U11036 ( .A1(n11123), .A2(n11124), .Y(n11122) );
  OR2X1_RVT U11037 ( .A1(n12226), .A2(n124), .Y(n11124) );
  NAND2X1_RVT U11038 ( .A1(n10609), .A2(n12839), .Y(n11123) );
  OR2X1_RVT U11039 ( .A1(n11125), .A2(n116), .Y(n11120) );
  AND2X1_RVT U11040 ( .A1(n10833), .A2(n10710), .Y(n11125) );
  OR2X1_RVT U11041 ( .A1(n10559), .A2(n11126), .Y(n10710) );
  OR2X1_RVT U11042 ( .A1(n12850), .A2(n12215), .Y(n11126) );
  AND4X1_RVT U11043 ( .A1(n10727), .A2(n11127), .A3(n10919), .A4(n11128), .Y(
        n11091) );
  AND4X1_RVT U11044 ( .A1(n11129), .A2(n11130), .A3(n11131), .A4(n11132), .Y(
        n11128) );
  OR2X1_RVT U11045 ( .A1(n10690), .A2(n10611), .Y(n11132) );
  OR2X1_RVT U11046 ( .A1(n10628), .A2(n10657), .Y(n11131) );
  OR2X1_RVT U11047 ( .A1(n12838), .A2(n10882), .Y(n11130) );
  OR2X1_RVT U11048 ( .A1(n10606), .A2(n10588), .Y(n10882) );
  OR2X1_RVT U11049 ( .A1(n12846), .A2(n10670), .Y(n10588) );
  OR2X1_RVT U11050 ( .A1(n12229), .A2(n10711), .Y(n11129) );
  OR2X1_RVT U11051 ( .A1(n10592), .A2(n10820), .Y(n10711) );
  OR2X1_RVT U11052 ( .A1(n12213), .A2(n10796), .Y(n10820) );
  AND2X1_RVT U11053 ( .A1(n11133), .A2(n11134), .Y(n10919) );
  OR2X1_RVT U11054 ( .A1(n11135), .A2(n10659), .Y(n11134) );
  OR2X1_RVT U11055 ( .A1(n12239), .A2(n116), .Y(n11135) );
  OR2X1_RVT U11056 ( .A1(n11136), .A2(n10542), .Y(n11133) );
  OR2X1_RVT U11057 ( .A1(n12837), .A2(n10659), .Y(n10542) );
  OR2X1_RVT U11058 ( .A1(n10556), .A2(n10606), .Y(n11136) );
  OR2X1_RVT U11059 ( .A1(n12221), .A2(n10925), .Y(n11127) );
  AND2X1_RVT U11060 ( .A1(n11137), .A2(n11138), .Y(n10727) );
  OR2X1_RVT U11061 ( .A1(n10610), .A2(n10648), .Y(n11138) );
  OR2X1_RVT U11062 ( .A1(n11139), .A2(n11140), .Y(n11137) );
  AND4X1_RVT U11063 ( .A1(n11141), .A2(n11142), .A3(n11143), .A4(n11144), .Y(
        n11090) );
  OR2X1_RVT U11064 ( .A1(n11145), .A2(n10796), .Y(n11144) );
  AND2X1_RVT U11065 ( .A1(n11146), .A2(n10805), .Y(n11145) );
  OR2X1_RVT U11066 ( .A1(n12227), .A2(n11102), .Y(n10805) );
  OR2X1_RVT U11067 ( .A1(n11147), .A2(n12843), .Y(n11143) );
  AND2X1_RVT U11068 ( .A1(n10733), .A2(n10698), .Y(n11147) );
  OR2X1_RVT U11069 ( .A1(n12837), .A2(n10674), .Y(n10698) );
  OR2X1_RVT U11070 ( .A1(n11148), .A2(n10753), .Y(n11142) );
  AND2X1_RVT U11071 ( .A1(n11149), .A2(n11150), .Y(n11148) );
  OR2X1_RVT U11072 ( .A1(n12216), .A2(n10612), .Y(n11150) );
  AND2X1_RVT U11073 ( .A1(n11151), .A2(n10650), .Y(n11149) );
  OR2X1_RVT U11074 ( .A1(n114), .A2(n10609), .Y(n11151) );
  OR2X1_RVT U11075 ( .A1(n11152), .A2(n10550), .Y(n11141) );
  AND2X1_RVT U11076 ( .A1(n11153), .A2(n11154), .Y(n11152) );
  NAND2X1_RVT U11077 ( .A1(n10535), .A2(n10913), .Y(n11154) );
  AND2X1_RVT U11078 ( .A1(n11155), .A2(n10763), .Y(n11153) );
  OR2X1_RVT U11079 ( .A1(n10696), .A2(n11102), .Y(n10763) );
  OR2X1_RVT U11080 ( .A1(n12236), .A2(n11156), .Y(n11155) );
  AND4X1_RVT U11081 ( .A1(n11157), .A2(n11158), .A3(n11159), .A4(n11160), .Y(
        n11089) );
  OR2X1_RVT U11082 ( .A1(n11161), .A2(n10573), .Y(n11160) );
  AND2X1_RVT U11083 ( .A1(n11162), .A2(n10714), .Y(n11161) );
  AND2X1_RVT U11084 ( .A1(n11163), .A2(n10736), .Y(n11162) );
  OR2X1_RVT U11085 ( .A1(n116), .A2(n11140), .Y(n10736) );
  OR2X1_RVT U11086 ( .A1(n12215), .A2(n10670), .Y(n11140) );
  OR2X1_RVT U11087 ( .A1(n11164), .A2(n12232), .Y(n11159) );
  AND2X1_RVT U11088 ( .A1(n11165), .A2(n11166), .Y(n11164) );
  OR2X1_RVT U11089 ( .A1(n11167), .A2(n12835), .Y(n11166) );
  AND2X1_RVT U11090 ( .A1(n11168), .A2(n11169), .Y(n11167) );
  OR2X1_RVT U11091 ( .A1(n12214), .A2(n10947), .Y(n11169) );
  OR2X1_RVT U11092 ( .A1(n12842), .A2(n10593), .Y(n11168) );
  AND2X1_RVT U11093 ( .A1(n11170), .A2(n11171), .Y(n11165) );
  OR2X1_RVT U11094 ( .A1(n10559), .A2(n11172), .Y(n11170) );
  OR2X1_RVT U11095 ( .A1(n11173), .A2(n10593), .Y(n11158) );
  AND4X1_RVT U11096 ( .A1(n11174), .A2(n11175), .A3(n11176), .A4(n10559), .Y(
        n11173) );
  OR2X1_RVT U11097 ( .A1(n12843), .A2(n10609), .Y(n11176) );
  OR2X1_RVT U11098 ( .A1(n12226), .A2(n10628), .Y(n11175) );
  OR2X1_RVT U11099 ( .A1(n10681), .A2(n10659), .Y(n11174) );
  OR2X1_RVT U11100 ( .A1(n11177), .A2(n10535), .Y(n11157) );
  AND4X1_RVT U11101 ( .A1(n10960), .A2(n11178), .A3(n10758), .A4(n10674), .Y(
        n11177) );
  OR2X1_RVT U11102 ( .A1(n10628), .A2(n11172), .Y(n10758) );
  OR2X1_RVT U11103 ( .A1(n10796), .A2(n11003), .Y(n11178) );
  OR2X1_RVT U11104 ( .A1(n12220), .A2(n10761), .Y(n10960) );
  AND4X1_RVT U11105 ( .A1(n11180), .A2(n11181), .A3(n11182), .A4(n11183), .Y(
        n11179) );
  AND4X1_RVT U11106 ( .A1(n10611), .A2(n10847), .A3(n11184), .A4(n11185), .Y(
        n11183) );
  AND4X1_RVT U11107 ( .A1(n10926), .A2(n10871), .A3(n11097), .A4(n11098), .Y(
        n11185) );
  OR2X1_RVT U11108 ( .A1(n11100), .A2(n10532), .Y(n11098) );
  OR2X1_RVT U11109 ( .A1(n12841), .A2(n10650), .Y(n10532) );
  OR2X1_RVT U11110 ( .A1(n10549), .A2(n11139), .Y(n11097) );
  OR2X1_RVT U11111 ( .A1(n12846), .A2(n12234), .Y(n11139) );
  OR2X1_RVT U11112 ( .A1(n12835), .A2(n10670), .Y(n10549) );
  OR2X1_RVT U11113 ( .A1(n12847), .A2(n10568), .Y(n10871) );
  OR2X1_RVT U11114 ( .A1(n12243), .A2(n12227), .Y(n10568) );
  OR2X1_RVT U11115 ( .A1(n10690), .A2(n11186), .Y(n10926) );
  OR2X1_RVT U11116 ( .A1(n12234), .A2(n10594), .Y(n11186) );
  OR2X1_RVT U11117 ( .A1(n10592), .A2(n11187), .Y(n11184) );
  OR2X1_RVT U11118 ( .A1(n10720), .A2(n12225), .Y(n11187) );
  OR2X1_RVT U11119 ( .A1(n10659), .A2(n11188), .Y(n10847) );
  OR2X1_RVT U11120 ( .A1(n10593), .A2(n12232), .Y(n11188) );
  OR2X1_RVT U11121 ( .A1(n12839), .A2(n11099), .Y(n10611) );
  OR2X1_RVT U11122 ( .A1(n12227), .A2(n10610), .Y(n11099) );
  AND4X1_RVT U11123 ( .A1(n11189), .A2(n11190), .A3(n11191), .A4(n11192), .Y(
        n11182) );
  AND4X1_RVT U11124 ( .A1(n11193), .A2(n11194), .A3(n11195), .A4(n11196), .Y(
        n11192) );
  OR2X1_RVT U11125 ( .A1(n10626), .A2(n11197), .Y(n11196) );
  OR2X1_RVT U11126 ( .A1(n12216), .A2(n10696), .Y(n11197) );
  OR2X1_RVT U11127 ( .A1(n10609), .A2(n11198), .Y(n11195) );
  OR2X1_RVT U11128 ( .A1(n11199), .A2(n10573), .Y(n11198) );
  AND2X1_RVT U11129 ( .A1(n10552), .A2(n10612), .Y(n11199) );
  OR2X1_RVT U11130 ( .A1(n11200), .A2(n11201), .Y(n11194) );
  AND2X1_RVT U11131 ( .A1(n10767), .A2(n10723), .Y(n11200) );
  OR2X1_RVT U11132 ( .A1(n12840), .A2(n124), .Y(n10723) );
  OR2X1_RVT U11133 ( .A1(n12836), .A2(n12237), .Y(n10767) );
  OR2X1_RVT U11134 ( .A1(n11202), .A2(n10607), .Y(n11193) );
  AND2X1_RVT U11135 ( .A1(n11003), .A2(n11203), .Y(n11202) );
  OR2X1_RVT U11136 ( .A1(n12838), .A2(n116), .Y(n11203) );
  OR2X1_RVT U11137 ( .A1(n11204), .A2(n12239), .Y(n11191) );
  AND2X1_RVT U11138 ( .A1(n10994), .A2(n11205), .Y(n11204) );
  OR2X1_RVT U11139 ( .A1(n10600), .A2(n10947), .Y(n11205) );
  OR2X1_RVT U11140 ( .A1(n12220), .A2(n10812), .Y(n10994) );
  OR2X1_RVT U11141 ( .A1(n12842), .A2(n10600), .Y(n10812) );
  OR2X1_RVT U11142 ( .A1(n11206), .A2(n10761), .Y(n11190) );
  AND2X1_RVT U11143 ( .A1(n10714), .A2(n10986), .Y(n11206) );
  OR2X1_RVT U11144 ( .A1(n10570), .A2(n10659), .Y(n10714) );
  OR2X1_RVT U11145 ( .A1(n11207), .A2(n10650), .Y(n11189) );
  AND2X1_RVT U11146 ( .A1(n10613), .A2(n10615), .Y(n11207) );
  AND4X1_RVT U11147 ( .A1(n11208), .A2(n11209), .A3(n11210), .A4(n11211), .Y(
        n11181) );
  AND4X1_RVT U11148 ( .A1(n11212), .A2(n11213), .A3(n11214), .A4(n11215), .Y(
        n11211) );
  OR2X1_RVT U11149 ( .A1(n11216), .A2(n12223), .Y(n11215) );
  AND2X1_RVT U11150 ( .A1(n10541), .A2(n10833), .Y(n11216) );
  OR2X1_RVT U11151 ( .A1(n10690), .A2(n10721), .Y(n10833) );
  OR2X1_RVT U11152 ( .A1(n12226), .A2(n10573), .Y(n10721) );
  OR2X1_RVT U11153 ( .A1(n12230), .A2(n11217), .Y(n10541) );
  OR2X1_RVT U11154 ( .A1(n12213), .A2(n12219), .Y(n11217) );
  OR2X1_RVT U11155 ( .A1(n11218), .A2(n12237), .Y(n11214) );
  AND2X1_RVT U11156 ( .A1(n10850), .A2(n11219), .Y(n11218) );
  OR2X1_RVT U11157 ( .A1(n12242), .A2(n114), .Y(n11219) );
  OR2X1_RVT U11158 ( .A1(n12240), .A2(n10657), .Y(n10850) );
  OR2X1_RVT U11159 ( .A1(n11220), .A2(n12218), .Y(n11213) );
  AND2X1_RVT U11160 ( .A1(n10868), .A2(n11221), .Y(n11220) );
  OR2X1_RVT U11161 ( .A1(n12243), .A2(n10593), .Y(n11221) );
  OR2X1_RVT U11162 ( .A1(n10535), .A2(n11222), .Y(n10868) );
  OR2X1_RVT U11163 ( .A1(n11223), .A2(n10594), .Y(n11212) );
  AND2X1_RVT U11164 ( .A1(n11224), .A2(n11225), .Y(n11223) );
  OR2X1_RVT U11165 ( .A1(n10650), .A2(n12240), .Y(n11225) );
  AND2X1_RVT U11166 ( .A1(n11226), .A2(n10626), .Y(n11224) );
  OR2X1_RVT U11167 ( .A1(n10612), .A2(n10573), .Y(n10626) );
  OR2X1_RVT U11168 ( .A1(n12215), .A2(n10657), .Y(n11226) );
  OR2X1_RVT U11169 ( .A1(n12850), .A2(n10612), .Y(n10657) );
  OR2X1_RVT U11170 ( .A1(n11227), .A2(n10670), .Y(n11210) );
  AND4X1_RVT U11171 ( .A1(n11228), .A2(n11229), .A3(n10823), .A4(n10733), .Y(
        n11227) );
  OR2X1_RVT U11172 ( .A1(n10796), .A2(n10896), .Y(n10733) );
  OR2X1_RVT U11173 ( .A1(n10628), .A2(n11156), .Y(n10823) );
  OR2X1_RVT U11174 ( .A1(n12221), .A2(n12214), .Y(n11156) );
  OR2X1_RVT U11175 ( .A1(n116), .A2(n10550), .Y(n11229) );
  OR2X1_RVT U11176 ( .A1(n114), .A2(n12240), .Y(n11228) );
  OR2X1_RVT U11177 ( .A1(n11230), .A2(n10606), .Y(n11209) );
  AND2X1_RVT U11178 ( .A1(n11231), .A2(n10627), .Y(n11230) );
  AND2X1_RVT U11179 ( .A1(n11163), .A2(n10877), .Y(n11231) );
  OR2X1_RVT U11180 ( .A1(n11232), .A2(n12847), .Y(n10877) );
  AND2X1_RVT U11181 ( .A1(n10648), .A2(n11233), .Y(n11232) );
  OR2X1_RVT U11182 ( .A1(n12218), .A2(n10535), .Y(n11233) );
  OR2X1_RVT U11183 ( .A1(n10696), .A2(n10834), .Y(n11163) );
  OR2X1_RVT U11184 ( .A1(n10681), .A2(n10570), .Y(n10834) );
  OR2X1_RVT U11185 ( .A1(n11234), .A2(n10674), .Y(n11208) );
  AND2X1_RVT U11186 ( .A1(n11235), .A2(n12226), .Y(n11234) );
  AND2X1_RVT U11187 ( .A1(n11236), .A2(n10855), .Y(n11235) );
  OR2X1_RVT U11188 ( .A1(n10696), .A2(n10796), .Y(n11236) );
  AND4X1_RVT U11189 ( .A1(n11237), .A2(n11238), .A3(n11239), .A4(n11240), .Y(
        n11180) );
  AND2X1_RVT U11190 ( .A1(n11241), .A2(n11242), .Y(n11240) );
  OR2X1_RVT U11191 ( .A1(n12843), .A2(n10776), .Y(n11242) );
  OR2X1_RVT U11192 ( .A1(n12234), .A2(n11243), .Y(n10776) );
  OR2X1_RVT U11193 ( .A1(n10592), .A2(n10681), .Y(n11243) );
  AND2X1_RVT U11194 ( .A1(n11244), .A2(n11245), .Y(n11241) );
  OR2X1_RVT U11195 ( .A1(n10565), .A2(n10576), .Y(n11245) );
  OR2X1_RVT U11196 ( .A1(n10609), .A2(n10804), .Y(n10576) );
  OR2X1_RVT U11197 ( .A1(n12839), .A2(n10570), .Y(n10804) );
  OR2X1_RVT U11198 ( .A1(n10612), .A2(n10689), .Y(n11244) );
  OR2X1_RVT U11199 ( .A1(n10600), .A2(n11246), .Y(n10689) );
  OR2X1_RVT U11200 ( .A1(n10600), .A2(n10780), .Y(n11239) );
  OR2X1_RVT U11201 ( .A1(n116), .A2(n12236), .Y(n10780) );
  OR2X1_RVT U11202 ( .A1(n11247), .A2(n10556), .Y(n11238) );
  AND4X1_RVT U11203 ( .A1(n11248), .A2(n11249), .A3(n11250), .A4(n11251), .Y(
        n11247) );
  OR2X1_RVT U11204 ( .A1(n12837), .A2(n11252), .Y(n11250) );
  OR2X1_RVT U11205 ( .A1(n11253), .A2(n12844), .Y(n11252) );
  AND2X1_RVT U11206 ( .A1(n10607), .A2(n11254), .Y(n11253) );
  OR2X1_RVT U11207 ( .A1(n12229), .A2(n11255), .Y(n11249) );
  OR2X1_RVT U11208 ( .A1(n10913), .A2(n10550), .Y(n11255) );
  OR2X1_RVT U11209 ( .A1(n10533), .A2(n10559), .Y(n11248) );
  OR2X1_RVT U11210 ( .A1(n12841), .A2(n10659), .Y(n10559) );
  OR2X1_RVT U11211 ( .A1(n11114), .A2(n10947), .Y(n11237) );
  OR2X1_RVT U11212 ( .A1(n12245), .A2(n10570), .Y(n10947) );
  AND4X1_RVT U11213 ( .A1(n11257), .A2(n11258), .A3(n11259), .A4(n11260), .Y(
        n11256) );
  AND4X1_RVT U11214 ( .A1(n11261), .A2(n11262), .A3(n11263), .A4(n11264), .Y(
        n11260) );
  AND4X1_RVT U11215 ( .A1(n11265), .A2(n11266), .A3(n11267), .A4(n11268), .Y(
        n11264) );
  OR2X1_RVT U11216 ( .A1(n11102), .A2(n11246), .Y(n11268) );
  OR2X1_RVT U11217 ( .A1(n12840), .A2(n12239), .Y(n11246) );
  OR2X1_RVT U11218 ( .A1(n12213), .A2(n12223), .Y(n11102) );
  OR2X1_RVT U11219 ( .A1(n11269), .A2(n10607), .Y(n11267) );
  AND2X1_RVT U11220 ( .A1(n10553), .A2(n11201), .Y(n11269) );
  OR2X1_RVT U11221 ( .A1(n116), .A2(n11270), .Y(n10553) );
  OR2X1_RVT U11222 ( .A1(n12213), .A2(n12837), .Y(n11270) );
  OR2X1_RVT U11223 ( .A1(n11271), .A2(n10535), .Y(n11266) );
  OR2X1_RVT U11224 ( .A1(n12227), .A2(n10696), .Y(n10535) );
  AND2X1_RVT U11225 ( .A1(n10671), .A2(n11272), .Y(n11271) );
  OR2X1_RVT U11226 ( .A1(n10550), .A2(n10752), .Y(n11272) );
  OR2X1_RVT U11227 ( .A1(n12231), .A2(n12219), .Y(n10550) );
  OR2X1_RVT U11228 ( .A1(n10796), .A2(n11273), .Y(n10671) );
  OR2X1_RVT U11229 ( .A1(n12848), .A2(n12234), .Y(n11273) );
  OR2X1_RVT U11230 ( .A1(n11274), .A2(n10594), .Y(n11265) );
  AND2X1_RVT U11231 ( .A1(n10991), .A2(n11275), .Y(n11274) );
  OR2X1_RVT U11232 ( .A1(n11276), .A2(n12837), .Y(n11275) );
  AND2X1_RVT U11233 ( .A1(n10650), .A2(n11003), .Y(n11276) );
  OR2X1_RVT U11234 ( .A1(n12845), .A2(n10612), .Y(n11003) );
  OR2X1_RVT U11235 ( .A1(n12240), .A2(n11277), .Y(n10991) );
  OR2X1_RVT U11236 ( .A1(n12850), .A2(n12846), .Y(n11277) );
  OR2X1_RVT U11237 ( .A1(n11278), .A2(n12218), .Y(n11263) );
  AND2X1_RVT U11238 ( .A1(n11279), .A2(n11280), .Y(n11278) );
  OR2X1_RVT U11239 ( .A1(n11281), .A2(n10696), .Y(n11280) );
  AND2X1_RVT U11240 ( .A1(n10761), .A2(n11282), .Y(n11281) );
  OR2X1_RVT U11241 ( .A1(n10552), .A2(n10674), .Y(n11279) );
  OR2X1_RVT U11242 ( .A1(n12232), .A2(n10610), .Y(n10674) );
  OR2X1_RVT U11243 ( .A1(n11283), .A2(n12846), .Y(n11262) );
  AND2X1_RVT U11244 ( .A1(n10766), .A2(n10925), .Y(n11283) );
  OR2X1_RVT U11245 ( .A1(n12230), .A2(n11284), .Y(n10925) );
  OR2X1_RVT U11246 ( .A1(n10606), .A2(n12219), .Y(n11284) );
  OR2X1_RVT U11247 ( .A1(n10552), .A2(n11114), .Y(n10766) );
  OR2X1_RVT U11248 ( .A1(n12219), .A2(n12234), .Y(n11114) );
  OR2X1_RVT U11249 ( .A1(n11285), .A2(n12216), .Y(n11261) );
  AND2X1_RVT U11250 ( .A1(n10806), .A2(n11286), .Y(n11285) );
  OR2X1_RVT U11251 ( .A1(n11101), .A2(n10600), .Y(n11286) );
  OR2X1_RVT U11252 ( .A1(n10659), .A2(n11222), .Y(n10806) );
  OR2X1_RVT U11253 ( .A1(n12845), .A2(n116), .Y(n11222) );
  AND2X1_RVT U11254 ( .A1(n12220), .A2(n12848), .Y(n10902) );
  AND4X1_RVT U11255 ( .A1(n11287), .A2(n11288), .A3(n11289), .A4(n11290), .Y(
        n11259) );
  AND4X1_RVT U11256 ( .A1(n11291), .A2(n11292), .A3(n11293), .A4(n11294), .Y(
        n11290) );
  OR2X1_RVT U11257 ( .A1(n11295), .A2(n12225), .Y(n11294) );
  AND2X1_RVT U11258 ( .A1(n10793), .A2(n10864), .Y(n11295) );
  OR2X1_RVT U11259 ( .A1(n10609), .A2(n11201), .Y(n10864) );
  OR2X1_RVT U11260 ( .A1(n12848), .A2(n10606), .Y(n11201) );
  OR2X1_RVT U11261 ( .A1(n12835), .A2(n12215), .Y(n10609) );
  OR2X1_RVT U11262 ( .A1(n12216), .A2(n10896), .Y(n10793) );
  OR2X1_RVT U11263 ( .A1(n12220), .A2(n12234), .Y(n10896) );
  OR2X1_RVT U11264 ( .A1(n11296), .A2(n12844), .Y(n11293) );
  AND2X1_RVT U11265 ( .A1(n10955), .A2(n11297), .Y(n11296) );
  OR2X1_RVT U11266 ( .A1(n10913), .A2(n10623), .Y(n11297) );
  OR2X1_RVT U11267 ( .A1(n10796), .A2(n11298), .Y(n10623) );
  OR2X1_RVT U11268 ( .A1(n12245), .A2(n12221), .Y(n11298) );
  OR2X1_RVT U11269 ( .A1(n12229), .A2(n11299), .Y(n10955) );
  OR2X1_RVT U11270 ( .A1(n10796), .A2(n10592), .Y(n11299) );
  OR2X1_RVT U11271 ( .A1(n11300), .A2(n12850), .Y(n11292) );
  AND2X1_RVT U11272 ( .A1(n10901), .A2(n10830), .Y(n11300) );
  OR2X1_RVT U11273 ( .A1(n10612), .A2(n10648), .Y(n10830) );
  OR2X1_RVT U11274 ( .A1(n12842), .A2(n10796), .Y(n10648) );
  OR2X1_RVT U11275 ( .A1(n11101), .A2(n10628), .Y(n10901) );
  OR2X1_RVT U11276 ( .A1(n12226), .A2(n12847), .Y(n11101) );
  OR2X1_RVT U11277 ( .A1(n11301), .A2(n10670), .Y(n11291) );
  AND2X1_RVT U11278 ( .A1(n11302), .A2(n11303), .Y(n11301) );
  OR2X1_RVT U11279 ( .A1(n10592), .A2(n11100), .Y(n11303) );
  OR2X1_RVT U11280 ( .A1(n12844), .A2(n124), .Y(n11100) );
  AND2X1_RVT U11281 ( .A1(n11304), .A2(n10887), .Y(n11302) );
  OR2X1_RVT U11282 ( .A1(n10600), .A2(n11305), .Y(n10887) );
  OR2X1_RVT U11283 ( .A1(n12242), .A2(n12221), .Y(n11305) );
  OR2X1_RVT U11284 ( .A1(n10656), .A2(n10593), .Y(n11289) );
  OR2X1_RVT U11285 ( .A1(n12837), .A2(n10552), .Y(n10656) );
  OR2X1_RVT U11286 ( .A1(n11306), .A2(n10556), .Y(n11288) );
  AND2X1_RVT U11287 ( .A1(n11307), .A2(n10737), .Y(n11306) );
  AND2X1_RVT U11288 ( .A1(n11308), .A2(n11309), .Y(n10737) );
  OR2X1_RVT U11289 ( .A1(n12230), .A2(n10761), .Y(n11309) );
  OR2X1_RVT U11290 ( .A1(n10659), .A2(n10533), .Y(n11308) );
  OR2X1_RVT U11291 ( .A1(n12215), .A2(n10606), .Y(n10533) );
  AND2X1_RVT U11292 ( .A1(n11310), .A2(n10923), .Y(n11307) );
  OR2X1_RVT U11293 ( .A1(n10690), .A2(n11254), .Y(n10923) );
  OR2X1_RVT U11294 ( .A1(n12839), .A2(n114), .Y(n11254) );
  OR2X1_RVT U11295 ( .A1(n10552), .A2(n10719), .Y(n11310) );
  OR2X1_RVT U11296 ( .A1(n12214), .A2(n11311), .Y(n10719) );
  OR2X1_RVT U11297 ( .A1(n12835), .A2(n12243), .Y(n11311) );
  OR2X1_RVT U11298 ( .A1(n11312), .A2(n12835), .Y(n11287) );
  AND4X1_RVT U11299 ( .A1(n11313), .A2(n11314), .A3(n11315), .A4(n11146), .Y(
        n11312) );
  OR2X1_RVT U11300 ( .A1(n10606), .A2(n10986), .Y(n11146) );
  OR2X1_RVT U11301 ( .A1(n12840), .A2(n12846), .Y(n10986) );
  OR2X1_RVT U11302 ( .A1(n10606), .A2(n11316), .Y(n11315) );
  OR2X1_RVT U11303 ( .A1(n12220), .A2(n12225), .Y(n11316) );
  OR2X1_RVT U11304 ( .A1(n12845), .A2(n10565), .Y(n10606) );
  OR2X1_RVT U11305 ( .A1(n11317), .A2(n10687), .Y(n11314) );
  OR2X1_RVT U11306 ( .A1(n12214), .A2(n10531), .Y(n10687) );
  AND2X1_RVT U11307 ( .A1(n10670), .A2(n11318), .Y(n11317) );
  OR2X1_RVT U11308 ( .A1(n12843), .A2(n10570), .Y(n11318) );
  OR2X1_RVT U11309 ( .A1(n12839), .A2(n12225), .Y(n10670) );
  OR2X1_RVT U11310 ( .A1(n12841), .A2(n11282), .Y(n11313) );
  OR2X1_RVT U11311 ( .A1(n12845), .A2(n10610), .Y(n11282) );
  OR2X1_RVT U11312 ( .A1(n10556), .A2(n114), .Y(n10610) );
  AND4X1_RVT U11313 ( .A1(n11319), .A2(n11320), .A3(n11321), .A4(n11322), .Y(
        n11258) );
  AND4X1_RVT U11314 ( .A1(n11323), .A2(n11324), .A3(n11325), .A4(n11326), .Y(
        n11322) );
  OR2X1_RVT U11315 ( .A1(n10628), .A2(n10755), .Y(n11326) );
  OR2X1_RVT U11316 ( .A1(n12227), .A2(n10650), .Y(n10755) );
  OR2X1_RVT U11317 ( .A1(n12231), .A2(n10796), .Y(n10628) );
  OR2X1_RVT U11318 ( .A1(n10615), .A2(n11172), .Y(n11325) );
  OR2X1_RVT U11319 ( .A1(n12849), .A2(n12214), .Y(n11172) );
  OR2X1_RVT U11320 ( .A1(n10681), .A2(n10607), .Y(n10615) );
  OR2X1_RVT U11321 ( .A1(n10600), .A2(n10627), .Y(n11324) );
  OR2X1_RVT U11322 ( .A1(n12223), .A2(n12236), .Y(n10627) );
  OR2X1_RVT U11323 ( .A1(n12213), .A2(n12836), .Y(n10600) );
  OR2X1_RVT U11324 ( .A1(n124), .A2(n10966), .Y(n11323) );
  OR2X1_RVT U11325 ( .A1(n12221), .A2(n10753), .Y(n10966) );
  OR2X1_RVT U11326 ( .A1(n10570), .A2(n11000), .Y(n11321) );
  OR2X1_RVT U11327 ( .A1(n124), .A2(n11327), .Y(n11000) );
  OR2X1_RVT U11328 ( .A1(n12842), .A2(n12234), .Y(n11327) );
  AND2X1_RVT U11329 ( .A1(n12215), .A2(n12218), .Y(n11111) );
  OR2X1_RVT U11330 ( .A1(n10612), .A2(n10560), .Y(n11320) );
  OR2X1_RVT U11331 ( .A1(n12243), .A2(n11328), .Y(n10560) );
  OR2X1_RVT U11332 ( .A1(n12843), .A2(n12835), .Y(n11328) );
  OR2X1_RVT U11333 ( .A1(n12220), .A2(n10592), .Y(n10612) );
  OR2X1_RVT U11334 ( .A1(n10659), .A2(n11304), .Y(n11319) );
  OR2X1_RVT U11335 ( .A1(n12216), .A2(n10614), .Y(n11304) );
  OR2X1_RVT U11336 ( .A1(n12845), .A2(n12846), .Y(n10614) );
  AND4X1_RVT U11337 ( .A1(n11329), .A2(n10725), .A3(n11330), .A4(n11331), .Y(
        n11257) );
  OR2X1_RVT U11338 ( .A1(n12220), .A2(n11251), .Y(n11331) );
  OR2X1_RVT U11339 ( .A1(n12841), .A2(n10720), .Y(n11251) );
  OR2X1_RVT U11340 ( .A1(n12218), .A2(n10761), .Y(n10720) );
  OR2X1_RVT U11341 ( .A1(n12213), .A2(n10587), .Y(n10761) );
  AND2X1_RVT U11342 ( .A1(n11332), .A2(n11333), .Y(n11330) );
  OR2X1_RVT U11343 ( .A1(n12242), .A2(n11171), .Y(n11333) );
  OR2X1_RVT U11344 ( .A1(n10659), .A2(n10752), .Y(n11171) );
  OR2X1_RVT U11345 ( .A1(n12220), .A2(n12214), .Y(n10752) );
  OR2X1_RVT U11346 ( .A1(n12215), .A2(n10548), .Y(n10587) );
  OR2X1_RVT U11347 ( .A1(n12848), .A2(n10821), .Y(n11332) );
  OR2X1_RVT U11348 ( .A1(n12239), .A2(n10855), .Y(n10821) );
  OR2X1_RVT U11349 ( .A1(n12840), .A2(n12835), .Y(n10855) );
  OR2X1_RVT U11350 ( .A1(n12838), .A2(n12231), .Y(n10531) );
  AND2X1_RVT U11351 ( .A1(n11334), .A2(n11335), .Y(n10725) );
  OR2X1_RVT U11352 ( .A1(n10607), .A2(n10593), .Y(n11335) );
  OR2X1_RVT U11353 ( .A1(n12847), .A2(n10565), .Y(n10593) );
  AND2X1_RVT U11354 ( .A1(n10592), .A2(n10556), .Y(n10645) );
  OR2X1_RVT U11355 ( .A1(n12226), .A2(n10659), .Y(n10607) );
  OR2X1_RVT U11356 ( .A1(n12836), .A2(n10696), .Y(n10659) );
  OR2X1_RVT U11357 ( .A1(n11336), .A2(n10650), .Y(n11334) );
  OR2X1_RVT U11358 ( .A1(n12220), .A2(n114), .Y(n10650) );
  AND2X1_RVT U11359 ( .A1(n12849), .A2(n12213), .Y(n10913) );
  OR2X1_RVT U11360 ( .A1(n12219), .A2(n10753), .Y(n11336) );
  OR2X1_RVT U11361 ( .A1(n12845), .A2(n12236), .Y(n10753) );
  AND2X1_RVT U11362 ( .A1(n11337), .A2(n11338), .Y(n11329) );
  OR2X1_RVT U11363 ( .A1(n10573), .A2(n10906), .Y(n11338) );
  OR2X1_RVT U11364 ( .A1(n12221), .A2(n10613), .Y(n10906) );
  OR2X1_RVT U11365 ( .A1(n12236), .A2(n10690), .Y(n10613) );
  OR2X1_RVT U11366 ( .A1(n12216), .A2(n12219), .Y(n10690) );
  OR2X1_RVT U11367 ( .A1(n12842), .A2(n12840), .Y(n10552) );
  OR2X1_RVT U11368 ( .A1(n12850), .A2(n12844), .Y(n10573) );
  XOR2X1_RVT U11369 ( .A1(key[84]), .A2(state[84]), .Y(n10548) );
  OR2X1_RVT U11370 ( .A1(n10565), .A2(n10694), .Y(n11337) );
  OR2X1_RVT U11371 ( .A1(n10796), .A2(n10987), .Y(n10694) );
  OR2X1_RVT U11372 ( .A1(n12223), .A2(n10594), .Y(n10987) );
  OR2X1_RVT U11373 ( .A1(n12843), .A2(n10696), .Y(n10594) );
  XOR2X1_RVT U11374 ( .A1(key[82]), .A2(state[82]), .Y(n10696) );
  XOR2X1_RVT U11375 ( .A1(key[83]), .A2(state[83]), .Y(n10630) );
  OR2X1_RVT U11376 ( .A1(n12848), .A2(n12221), .Y(n10570) );
  XOR2X1_RVT U11377 ( .A1(key[85]), .A2(state[85]), .Y(n10556) );
  XOR2X1_RVT U11378 ( .A1(key[86]), .A2(state[86]), .Y(n10592) );
  OR2X1_RVT U11379 ( .A1(n12838), .A2(n12219), .Y(n10796) );
  XOR2X1_RVT U11380 ( .A1(key[80]), .A2(state[80]), .Y(n10571) );
  XOR2X1_RVT U11381 ( .A1(key[81]), .A2(state[81]), .Y(n10681) );
  XOR2X1_RVT U11382 ( .A1(key[87]), .A2(state[87]), .Y(n10565) );
  AND4X1_RVT U11383 ( .A1(n11340), .A2(n11341), .A3(n11342), .A4(n11343), .Y(
        n11339) );
  AND4X1_RVT U11384 ( .A1(n11344), .A2(n11345), .A3(n11346), .A4(n11347), .Y(
        n11343) );
  AND4X1_RVT U11385 ( .A1(n11348), .A2(n11349), .A3(n11350), .A4(n11351), .Y(
        n11347) );
  OR2X1_RVT U11386 ( .A1(n12178), .A2(n11353), .Y(n11346) );
  OR2X1_RVT U11387 ( .A1(n11354), .A2(n11355), .Y(n11344) );
  OR2X1_RVT U11388 ( .A1(n12832), .A2(n11356), .Y(n11355) );
  AND4X1_RVT U11389 ( .A1(n11357), .A2(n11358), .A3(n11359), .A4(n11360), .Y(
        n11342) );
  OR2X1_RVT U11390 ( .A1(n11361), .A2(n12830), .Y(n11360) );
  AND2X1_RVT U11391 ( .A1(n11362), .A2(n11363), .Y(n11361) );
  AND2X1_RVT U11392 ( .A1(n11364), .A2(n11365), .Y(n11359) );
  OR2X1_RVT U11393 ( .A1(n11366), .A2(n136), .Y(n11365) );
  AND2X1_RVT U11394 ( .A1(n11367), .A2(n11368), .Y(n11366) );
  OR2X1_RVT U11395 ( .A1(n12169), .A2(n11370), .Y(n11368) );
  OR2X1_RVT U11396 ( .A1(n11356), .A2(n11371), .Y(n11367) );
  OR2X1_RVT U11397 ( .A1(n11372), .A2(n12175), .Y(n11364) );
  AND2X1_RVT U11398 ( .A1(n11374), .A2(n11375), .Y(n11372) );
  OR2X1_RVT U11399 ( .A1(n11376), .A2(n11377), .Y(n11358) );
  AND2X1_RVT U11400 ( .A1(n11378), .A2(n11379), .Y(n11376) );
  OR2X1_RVT U11401 ( .A1(n12170), .A2(n11380), .Y(n11379) );
  AND2X1_RVT U11402 ( .A1(n11381), .A2(n11382), .Y(n11378) );
  AND2X1_RVT U11403 ( .A1(n11383), .A2(n11384), .Y(n11357) );
  OR2X1_RVT U11404 ( .A1(n11385), .A2(n12152), .Y(n11384) );
  AND2X1_RVT U11405 ( .A1(n11387), .A2(n11388), .Y(n11385) );
  OR2X1_RVT U11406 ( .A1(n11389), .A2(n11390), .Y(n11388) );
  OR2X1_RVT U11407 ( .A1(n12161), .A2(n12156), .Y(n11390) );
  OR2X1_RVT U11408 ( .A1(n11393), .A2(n11394), .Y(n11383) );
  AND2X1_RVT U11409 ( .A1(n11395), .A2(n11396), .Y(n11393) );
  AND2X1_RVT U11410 ( .A1(n11397), .A2(n11398), .Y(n11395) );
  AND4X1_RVT U11411 ( .A1(n11399), .A2(n11400), .A3(n11401), .A4(n11402), .Y(
        n11341) );
  AND4X1_RVT U11412 ( .A1(n11403), .A2(n11404), .A3(n11405), .A4(n11406), .Y(
        n11402) );
  OR2X1_RVT U11413 ( .A1(n11407), .A2(n12181), .Y(n11406) );
  AND4X1_RVT U11414 ( .A1(n11409), .A2(n11410), .A3(n11411), .A4(n11412), .Y(
        n11407) );
  OR2X1_RVT U11415 ( .A1(n11413), .A2(n11380), .Y(n11412) );
  OR2X1_RVT U11416 ( .A1(n11414), .A2(n12167), .Y(n11411) );
  OR2X1_RVT U11417 ( .A1(n11416), .A2(n12158), .Y(n11405) );
  AND4X1_RVT U11418 ( .A1(n11417), .A2(n11418), .A3(n11419), .A4(n11420), .Y(
        n11416) );
  OR2X1_RVT U11419 ( .A1(n11421), .A2(n11422), .Y(n11420) );
  OR2X1_RVT U11420 ( .A1(n12175), .A2(n12170), .Y(n11422) );
  AND2X1_RVT U11421 ( .A1(n11423), .A2(n11424), .Y(n11419) );
  OR2X1_RVT U11422 ( .A1(n12834), .A2(n11425), .Y(n11418) );
  OR2X1_RVT U11423 ( .A1(n11426), .A2(n11427), .Y(n11417) );
  AND2X1_RVT U11424 ( .A1(n11428), .A2(n11429), .Y(n11426) );
  OR2X1_RVT U11425 ( .A1(n12175), .A2(n11430), .Y(n11429) );
  OR2X1_RVT U11426 ( .A1(n11363), .A2(n11431), .Y(n11404) );
  OR2X1_RVT U11427 ( .A1(n11430), .A2(n11432), .Y(n11403) );
  OR2X1_RVT U11428 ( .A1(n11433), .A2(n11434), .Y(n11401) );
  OR2X1_RVT U11429 ( .A1(n11435), .A2(n11428), .Y(n11400) );
  OR2X1_RVT U11430 ( .A1(n11436), .A2(n11437), .Y(n11399) );
  AND4X1_RVT U11431 ( .A1(n11438), .A2(n11439), .A3(n11440), .A4(n11441), .Y(
        n11340) );
  AND2X1_RVT U11432 ( .A1(n11442), .A2(n11443), .Y(n11441) );
  OR2X1_RVT U11433 ( .A1(n11427), .A2(n11444), .Y(n11443) );
  AND2X1_RVT U11434 ( .A1(n11445), .A2(n11446), .Y(n11442) );
  OR2X1_RVT U11435 ( .A1(n11447), .A2(n11370), .Y(n11446) );
  OR2X1_RVT U11436 ( .A1(n11371), .A2(n11448), .Y(n11445) );
  OR2X1_RVT U11437 ( .A1(n134), .A2(n11449), .Y(n11440) );
  OR2X1_RVT U11438 ( .A1(n11450), .A2(n12165), .Y(n11439) );
  OR2X1_RVT U11439 ( .A1(n12168), .A2(n11452), .Y(n11438) );
  AND4X1_RVT U11440 ( .A1(n11454), .A2(n11455), .A3(n11456), .A4(n11457), .Y(
        n11453) );
  AND4X1_RVT U11441 ( .A1(n11458), .A2(n11349), .A3(n11459), .A4(n11460), .Y(
        n11457) );
  AND4X1_RVT U11442 ( .A1(n11461), .A2(n11462), .A3(n11463), .A4(n11464), .Y(
        n11460) );
  OR2X1_RVT U11443 ( .A1(n11370), .A2(n11465), .Y(n11464) );
  OR2X1_RVT U11444 ( .A1(n11466), .A2(n12180), .Y(n11465) );
  OR2X1_RVT U11445 ( .A1(n11371), .A2(n11467), .Y(n11463) );
  OR2X1_RVT U11446 ( .A1(n134), .A2(n12164), .Y(n11467) );
  OR2X1_RVT U11447 ( .A1(n11468), .A2(n11414), .Y(n11462) );
  AND2X1_RVT U11448 ( .A1(n11425), .A2(n11469), .Y(n11468) );
  OR2X1_RVT U11449 ( .A1(n11470), .A2(n11471), .Y(n11461) );
  AND2X1_RVT U11450 ( .A1(n11472), .A2(n11473), .Y(n11470) );
  AND2X1_RVT U11451 ( .A1(n11474), .A2(n11475), .Y(n11459) );
  OR2X1_RVT U11452 ( .A1(n11421), .A2(n11476), .Y(n11475) );
  OR2X1_RVT U11453 ( .A1(n11477), .A2(n12832), .Y(n11476) );
  OR2X1_RVT U11454 ( .A1(n11478), .A2(n11479), .Y(n11474) );
  OR2X1_RVT U11455 ( .A1(n11480), .A2(n12169), .Y(n11479) );
  OR2X1_RVT U11456 ( .A1(n11356), .A2(n11481), .Y(n11349) );
  AND4X1_RVT U11457 ( .A1(n11482), .A2(n11483), .A3(n11484), .A4(n11485), .Y(
        n11456) );
  AND4X1_RVT U11458 ( .A1(n11486), .A2(n11487), .A3(n11488), .A4(n11489), .Y(
        n11485) );
  OR2X1_RVT U11459 ( .A1(n11490), .A2(n12183), .Y(n11489) );
  AND2X1_RVT U11460 ( .A1(n11492), .A2(n11493), .Y(n11490) );
  OR2X1_RVT U11461 ( .A1(n12152), .A2(n11371), .Y(n11493) );
  OR2X1_RVT U11462 ( .A1(n11494), .A2(n11373), .Y(n11488) );
  AND2X1_RVT U11463 ( .A1(n11495), .A2(n11496), .Y(n11494) );
  OR2X1_RVT U11464 ( .A1(n11497), .A2(n12831), .Y(n11487) );
  AND2X1_RVT U11465 ( .A1(n11498), .A2(n11499), .Y(n11497) );
  OR2X1_RVT U11466 ( .A1(n11500), .A2(n11449), .Y(n11499) );
  AND2X1_RVT U11467 ( .A1(n12183), .A2(n12167), .Y(n11500) );
  OR2X1_RVT U11468 ( .A1(n11501), .A2(n12153), .Y(n11486) );
  AND2X1_RVT U11469 ( .A1(n11503), .A2(n11504), .Y(n11501) );
  OR2X1_RVT U11470 ( .A1(n11505), .A2(n12159), .Y(n11484) );
  AND2X1_RVT U11471 ( .A1(n11506), .A2(n11507), .Y(n11505) );
  OR2X1_RVT U11472 ( .A1(n12167), .A2(n11508), .Y(n11507) );
  AND2X1_RVT U11473 ( .A1(n11509), .A2(n11510), .Y(n11506) );
  OR2X1_RVT U11474 ( .A1(n11511), .A2(n11512), .Y(n11509) );
  OR2X1_RVT U11475 ( .A1(n11356), .A2(n11427), .Y(n11512) );
  OR2X1_RVT U11476 ( .A1(n11513), .A2(n12828), .Y(n11483) );
  AND2X1_RVT U11477 ( .A1(n11514), .A2(n11515), .Y(n11513) );
  OR2X1_RVT U11478 ( .A1(n11516), .A2(n11517), .Y(n11482) );
  AND2X1_RVT U11479 ( .A1(n11518), .A2(n11519), .Y(n11516) );
  AND2X1_RVT U11480 ( .A1(n11520), .A2(n11521), .Y(n11518) );
  OR2X1_RVT U11481 ( .A1(n136), .A2(n11449), .Y(n11521) );
  OR2X1_RVT U11482 ( .A1(n12177), .A2(n11414), .Y(n11520) );
  AND4X1_RVT U11483 ( .A1(n11522), .A2(n11523), .A3(n11524), .A4(n11525), .Y(
        n11455) );
  AND4X1_RVT U11484 ( .A1(n11526), .A2(n11527), .A3(n11528), .A4(n11529), .Y(
        n11525) );
  OR2X1_RVT U11485 ( .A1(n11449), .A2(n11448), .Y(n11529) );
  OR2X1_RVT U11486 ( .A1(n11380), .A2(n11530), .Y(n11528) );
  OR2X1_RVT U11487 ( .A1(n11413), .A2(n11531), .Y(n11527) );
  OR2X1_RVT U11488 ( .A1(n11356), .A2(n11532), .Y(n11526) );
  AND2X1_RVT U11489 ( .A1(n11533), .A2(n11534), .Y(n11524) );
  OR2X1_RVT U11490 ( .A1(n12178), .A2(n11535), .Y(n11534) );
  OR2X1_RVT U11491 ( .A1(n12157), .A2(n11432), .Y(n11533) );
  OR2X1_RVT U11492 ( .A1(n11536), .A2(n11391), .Y(n11523) );
  AND4X1_RVT U11493 ( .A1(n11537), .A2(n11538), .A3(n11539), .A4(n11540), .Y(
        n11536) );
  OR2X1_RVT U11494 ( .A1(n11541), .A2(n11356), .Y(n11539) );
  OR2X1_RVT U11495 ( .A1(n12820), .A2(n11542), .Y(n11538) );
  OR2X1_RVT U11496 ( .A1(n11543), .A2(n12828), .Y(n11537) );
  AND2X1_RVT U11497 ( .A1(n11434), .A2(n11544), .Y(n11543) );
  OR2X1_RVT U11498 ( .A1(n11436), .A2(n11545), .Y(n11522) );
  AND4X1_RVT U11499 ( .A1(n11546), .A2(n11547), .A3(n11548), .A4(n11549), .Y(
        n11454) );
  AND4X1_RVT U11500 ( .A1(n11550), .A2(n11551), .A3(n11552), .A4(n11553), .Y(
        n11549) );
  OR2X1_RVT U11501 ( .A1(n12824), .A2(n11554), .Y(n11553) );
  OR2X1_RVT U11502 ( .A1(n12825), .A2(n11555), .Y(n11552) );
  OR2X1_RVT U11503 ( .A1(n12822), .A2(n11556), .Y(n11551) );
  OR2X1_RVT U11504 ( .A1(n12151), .A2(n11557), .Y(n11550) );
  OR2X1_RVT U11505 ( .A1(n11558), .A2(n12158), .Y(n11547) );
  AND4X1_RVT U11506 ( .A1(n11560), .A2(n11561), .A3(n11562), .A4(n11563), .Y(
        n11559) );
  AND4X1_RVT U11507 ( .A1(n11564), .A2(n11565), .A3(n11566), .A4(n11567), .Y(
        n11563) );
  AND4X1_RVT U11508 ( .A1(n11568), .A2(n11345), .A3(n11515), .A4(n11569), .Y(
        n11567) );
  OR2X1_RVT U11509 ( .A1(n11570), .A2(n12819), .Y(n11345) );
  AND2X1_RVT U11510 ( .A1(n11571), .A2(n11572), .Y(n11570) );
  OR2X1_RVT U11511 ( .A1(n11389), .A2(n11573), .Y(n11572) );
  OR2X1_RVT U11512 ( .A1(n11574), .A2(n11471), .Y(n11571) );
  OR2X1_RVT U11513 ( .A1(n11575), .A2(n11430), .Y(n11568) );
  AND2X1_RVT U11514 ( .A1(n11576), .A2(n11577), .Y(n11575) );
  OR2X1_RVT U11515 ( .A1(n12824), .A2(n11414), .Y(n11577) );
  OR2X1_RVT U11516 ( .A1(n11578), .A2(n11373), .Y(n11566) );
  AND2X1_RVT U11517 ( .A1(n11579), .A2(n11580), .Y(n11578) );
  OR2X1_RVT U11518 ( .A1(n11581), .A2(n12830), .Y(n11580) );
  AND2X1_RVT U11519 ( .A1(n11421), .A2(n11582), .Y(n11581) );
  OR2X1_RVT U11520 ( .A1(n11583), .A2(n12178), .Y(n11565) );
  AND2X1_RVT U11521 ( .A1(n11584), .A2(n11585), .Y(n11583) );
  OR2X1_RVT U11522 ( .A1(n11414), .A2(n11380), .Y(n11585) );
  OR2X1_RVT U11523 ( .A1(n11586), .A2(n12161), .Y(n11564) );
  AND2X1_RVT U11524 ( .A1(n11498), .A2(n11587), .Y(n11586) );
  OR2X1_RVT U11525 ( .A1(n11427), .A2(n11588), .Y(n11498) );
  AND4X1_RVT U11526 ( .A1(n11589), .A2(n11590), .A3(n11591), .A4(n11592), .Y(
        n11562) );
  OR2X1_RVT U11527 ( .A1(n11593), .A2(n12168), .Y(n11592) );
  AND2X1_RVT U11528 ( .A1(n11594), .A2(n11595), .Y(n11593) );
  OR2X1_RVT U11529 ( .A1(n11471), .A2(n11371), .Y(n11595) );
  AND2X1_RVT U11530 ( .A1(n11596), .A2(n11597), .Y(n11594) );
  OR2X1_RVT U11531 ( .A1(n11511), .A2(n11573), .Y(n11596) );
  AND2X1_RVT U11532 ( .A1(n11598), .A2(n11599), .Y(n11591) );
  OR2X1_RVT U11533 ( .A1(n11600), .A2(n11502), .Y(n11599) );
  AND2X1_RVT U11534 ( .A1(n11601), .A2(n11410), .Y(n11600) );
  OR2X1_RVT U11535 ( .A1(n11356), .A2(n11471), .Y(n11410) );
  OR2X1_RVT U11536 ( .A1(n11602), .A2(n136), .Y(n11598) );
  AND2X1_RVT U11537 ( .A1(n11603), .A2(n11604), .Y(n11602) );
  OR2X1_RVT U11538 ( .A1(n11605), .A2(n12170), .Y(n11604) );
  AND2X1_RVT U11539 ( .A1(n11606), .A2(n11607), .Y(n11605) );
  OR2X1_RVT U11540 ( .A1(n12165), .A2(n11421), .Y(n11607) );
  OR2X1_RVT U11541 ( .A1(n12834), .A2(n12167), .Y(n11606) );
  AND2X1_RVT U11542 ( .A1(n11472), .A2(n11582), .Y(n11603) );
  OR2X1_RVT U11543 ( .A1(n11502), .A2(n11608), .Y(n11472) );
  OR2X1_RVT U11544 ( .A1(n12829), .A2(n12825), .Y(n11608) );
  OR2X1_RVT U11545 ( .A1(n11609), .A2(n11491), .Y(n11590) );
  AND4X1_RVT U11546 ( .A1(n11450), .A2(n11610), .A3(n11611), .A4(n11612), .Y(
        n11609) );
  OR2X1_RVT U11547 ( .A1(n12169), .A2(n11471), .Y(n11612) );
  AND2X1_RVT U11548 ( .A1(n11613), .A2(n11614), .Y(n11611) );
  OR2X1_RVT U11549 ( .A1(n12834), .A2(n12178), .Y(n11610) );
  AND2X1_RVT U11550 ( .A1(n11615), .A2(n11616), .Y(n11450) );
  OR2X1_RVT U11551 ( .A1(n11617), .A2(n134), .Y(n11616) );
  OR2X1_RVT U11552 ( .A1(n11414), .A2(n12819), .Y(n11615) );
  AND2X1_RVT U11553 ( .A1(n11618), .A2(n11619), .Y(n11589) );
  OR2X1_RVT U11554 ( .A1(n11620), .A2(n12821), .Y(n11619) );
  AND2X1_RVT U11555 ( .A1(n11621), .A2(n11622), .Y(n11620) );
  OR2X1_RVT U11556 ( .A1(n11623), .A2(n12172), .Y(n11622) );
  AND2X1_RVT U11557 ( .A1(n11624), .A2(n11625), .Y(n11623) );
  AND2X1_RVT U11558 ( .A1(n11626), .A2(n11627), .Y(n11621) );
  OR2X1_RVT U11559 ( .A1(n11628), .A2(n12181), .Y(n11618) );
  AND4X1_RVT U11560 ( .A1(n11629), .A2(n11630), .A3(n11631), .A4(n11632), .Y(
        n11628) );
  OR2X1_RVT U11561 ( .A1(n12833), .A2(n11633), .Y(n11631) );
  OR2X1_RVT U11562 ( .A1(n134), .A2(n11428), .Y(n11630) );
  OR2X1_RVT U11563 ( .A1(n11517), .A2(n11471), .Y(n11629) );
  AND4X1_RVT U11564 ( .A1(n11634), .A2(n11635), .A3(n11636), .A4(n11637), .Y(
        n11561) );
  AND2X1_RVT U11565 ( .A1(n11638), .A2(n11481), .Y(n11637) );
  OR2X1_RVT U11566 ( .A1(n12156), .A2(n11447), .Y(n11481) );
  AND2X1_RVT U11567 ( .A1(n11639), .A2(n11640), .Y(n11638) );
  OR2X1_RVT U11568 ( .A1(n11641), .A2(n11396), .Y(n11640) );
  OR2X1_RVT U11569 ( .A1(n11448), .A2(n11508), .Y(n11639) );
  OR2X1_RVT U11570 ( .A1(n134), .A2(n11642), .Y(n11636) );
  OR2X1_RVT U11571 ( .A1(n12832), .A2(n11643), .Y(n11635) );
  OR2X1_RVT U11572 ( .A1(n11517), .A2(n11644), .Y(n11634) );
  AND4X1_RVT U11573 ( .A1(n11645), .A2(n11646), .A3(n11647), .A4(n11648), .Y(
        n11560) );
  AND2X1_RVT U11574 ( .A1(n11649), .A2(n11650), .Y(n11648) );
  OR2X1_RVT U11575 ( .A1(n12151), .A2(n11651), .Y(n11650) );
  AND2X1_RVT U11576 ( .A1(n11652), .A2(n11653), .Y(n11649) );
  OR2X1_RVT U11577 ( .A1(n11413), .A2(n11423), .Y(n11653) );
  OR2X1_RVT U11578 ( .A1(n12172), .A2(n11473), .Y(n11423) );
  OR2X1_RVT U11579 ( .A1(n12158), .A2(n11654), .Y(n11652) );
  OR2X1_RVT U11580 ( .A1(n11394), .A2(n11387), .Y(n11647) );
  OR2X1_RVT U11581 ( .A1(n11480), .A2(n11655), .Y(n11387) );
  OR2X1_RVT U11582 ( .A1(n12828), .A2(n11656), .Y(n11646) );
  OR2X1_RVT U11583 ( .A1(n12170), .A2(n11514), .Y(n11645) );
  OR2X1_RVT U11584 ( .A1(n12819), .A2(n11576), .Y(n11514) );
  AND4X1_RVT U11585 ( .A1(n11658), .A2(n11659), .A3(n11660), .A4(n11661), .Y(
        n11657) );
  AND4X1_RVT U11586 ( .A1(n11662), .A2(n11663), .A3(n11664), .A4(n11665), .Y(
        n11661) );
  OR2X1_RVT U11587 ( .A1(n144), .A2(n11666), .Y(n11665) );
  OR2X1_RVT U11588 ( .A1(n11667), .A2(n12183), .Y(n11666) );
  AND2X1_RVT U11589 ( .A1(n12172), .A2(n11433), .Y(n11667) );
  AND2X1_RVT U11590 ( .A1(n11348), .A2(n11668), .Y(n11664) );
  OR2X1_RVT U11591 ( .A1(n12161), .A2(n11669), .Y(n11348) );
  OR2X1_RVT U11592 ( .A1(n144), .A2(n11427), .Y(n11669) );
  OR2X1_RVT U11593 ( .A1(n11670), .A2(n11356), .Y(n11663) );
  AND2X1_RVT U11594 ( .A1(n11671), .A2(n11672), .Y(n11670) );
  AND2X1_RVT U11595 ( .A1(n11673), .A2(n11674), .Y(n11662) );
  OR2X1_RVT U11596 ( .A1(n11675), .A2(n11676), .Y(n11674) );
  AND2X1_RVT U11597 ( .A1(n11677), .A2(n11437), .Y(n11675) );
  OR2X1_RVT U11598 ( .A1(n11678), .A2(n11428), .Y(n11673) );
  AND2X1_RVT U11599 ( .A1(n11613), .A2(n11447), .Y(n11678) );
  OR2X1_RVT U11600 ( .A1(n12159), .A2(n11679), .Y(n11613) );
  OR2X1_RVT U11601 ( .A1(n12834), .A2(n12169), .Y(n11679) );
  AND4X1_RVT U11602 ( .A1(n11680), .A2(n11681), .A3(n11682), .A4(n11683), .Y(
        n11660) );
  OR2X1_RVT U11603 ( .A1(n11684), .A2(n12824), .Y(n11683) );
  AND2X1_RVT U11604 ( .A1(n11496), .A2(n11685), .Y(n11684) );
  OR2X1_RVT U11605 ( .A1(n12832), .A2(n11541), .Y(n11496) );
  AND2X1_RVT U11606 ( .A1(n11686), .A2(n11687), .Y(n11682) );
  OR2X1_RVT U11607 ( .A1(n11688), .A2(n12822), .Y(n11687) );
  AND2X1_RVT U11608 ( .A1(n11689), .A2(n11690), .Y(n11688) );
  OR2X1_RVT U11609 ( .A1(n11391), .A2(n11633), .Y(n11690) );
  OR2X1_RVT U11610 ( .A1(n11691), .A2(n12820), .Y(n11686) );
  AND2X1_RVT U11611 ( .A1(n11692), .A2(n11693), .Y(n11691) );
  OR2X1_RVT U11612 ( .A1(n11694), .A2(n12172), .Y(n11681) );
  AND2X1_RVT U11613 ( .A1(n11695), .A2(n11696), .Y(n11694) );
  AND2X1_RVT U11614 ( .A1(n11697), .A2(n11698), .Y(n11695) );
  AND2X1_RVT U11615 ( .A1(n11699), .A2(n11700), .Y(n11680) );
  OR2X1_RVT U11616 ( .A1(n11701), .A2(n11617), .Y(n11700) );
  AND2X1_RVT U11617 ( .A1(n11702), .A2(n11448), .Y(n11701) );
  AND2X1_RVT U11618 ( .A1(n11703), .A2(n11704), .Y(n11702) );
  OR2X1_RVT U11619 ( .A1(n11705), .A2(n12175), .Y(n11699) );
  AND2X1_RVT U11620 ( .A1(n11706), .A2(n11707), .Y(n11705) );
  OR2X1_RVT U11621 ( .A1(n12831), .A2(n12177), .Y(n11707) );
  AND2X1_RVT U11622 ( .A1(n11437), .A2(n11708), .Y(n11706) );
  AND4X1_RVT U11623 ( .A1(n11709), .A2(n11710), .A3(n11711), .A4(n11712), .Y(
        n11659) );
  AND2X1_RVT U11624 ( .A1(n11713), .A2(n11714), .Y(n11712) );
  OR2X1_RVT U11625 ( .A1(n11430), .A2(n11504), .Y(n11714) );
  OR2X1_RVT U11626 ( .A1(n12826), .A2(n11437), .Y(n11504) );
  AND2X1_RVT U11627 ( .A1(n11715), .A2(n11716), .Y(n11713) );
  OR2X1_RVT U11628 ( .A1(n11582), .A2(n11396), .Y(n11716) );
  OR2X1_RVT U11629 ( .A1(n12833), .A2(n12168), .Y(n11396) );
  OR2X1_RVT U11630 ( .A1(n11480), .A2(n11530), .Y(n11715) );
  OR2X1_RVT U11631 ( .A1(n12821), .A2(n11717), .Y(n11530) );
  OR2X1_RVT U11632 ( .A1(n11718), .A2(n12151), .Y(n11711) );
  AND4X1_RVT U11633 ( .A1(n11719), .A2(n11720), .A3(n11721), .A4(n11722), .Y(
        n11718) );
  OR2X1_RVT U11634 ( .A1(n11655), .A2(n11428), .Y(n11721) );
  OR2X1_RVT U11635 ( .A1(n11723), .A2(n11425), .Y(n11720) );
  OR2X1_RVT U11636 ( .A1(n12830), .A2(n11380), .Y(n11719) );
  OR2X1_RVT U11637 ( .A1(n11724), .A2(n12152), .Y(n11710) );
  AND2X1_RVT U11638 ( .A1(n11725), .A2(n11726), .Y(n11724) );
  OR2X1_RVT U11639 ( .A1(n11655), .A2(n11380), .Y(n11726) );
  AND2X1_RVT U11640 ( .A1(n11727), .A2(n11656), .Y(n11725) );
  OR2X1_RVT U11641 ( .A1(n11428), .A2(n11728), .Y(n11656) );
  OR2X1_RVT U11642 ( .A1(n12821), .A2(n12833), .Y(n11728) );
  OR2X1_RVT U11643 ( .A1(n11729), .A2(n12159), .Y(n11709) );
  AND4X1_RVT U11644 ( .A1(n11730), .A2(n11643), .A3(n11452), .A4(n11424), .Y(
        n11729) );
  OR2X1_RVT U11645 ( .A1(n11449), .A2(n11731), .Y(n11424) );
  OR2X1_RVT U11646 ( .A1(n12823), .A2(n11386), .Y(n11731) );
  OR2X1_RVT U11647 ( .A1(n11511), .A2(n11545), .Y(n11452) );
  OR2X1_RVT U11648 ( .A1(n11430), .A2(n11732), .Y(n11643) );
  OR2X1_RVT U11649 ( .A1(n12183), .A2(n12152), .Y(n11732) );
  OR2X1_RVT U11650 ( .A1(n11389), .A2(n11733), .Y(n11730) );
  OR2X1_RVT U11651 ( .A1(n11734), .A2(n12157), .Y(n11733) );
  AND4X1_RVT U11652 ( .A1(n11735), .A2(n11736), .A3(n11737), .A4(n11738), .Y(
        n11658) );
  AND2X1_RVT U11653 ( .A1(n11739), .A2(n11740), .Y(n11738) );
  AND2X1_RVT U11654 ( .A1(n11741), .A2(n11742), .Y(n11739) );
  OR2X1_RVT U11655 ( .A1(n11421), .A2(n11696), .Y(n11742) );
  OR2X1_RVT U11656 ( .A1(n11433), .A2(n11743), .Y(n11696) );
  OR2X1_RVT U11657 ( .A1(n12822), .A2(n12824), .Y(n11743) );
  OR2X1_RVT U11658 ( .A1(n12829), .A2(n11744), .Y(n11741) );
  OR2X1_RVT U11659 ( .A1(n12168), .A2(n11745), .Y(n11737) );
  OR2X1_RVT U11660 ( .A1(n12832), .A2(n11746), .Y(n11736) );
  OR2X1_RVT U11661 ( .A1(n11433), .A2(n11747), .Y(n11735) );
  AND4X1_RVT U11662 ( .A1(n11749), .A2(n11750), .A3(n11751), .A4(n11752), .Y(
        n11748) );
  AND4X1_RVT U11663 ( .A1(n11753), .A2(n11754), .A3(n11755), .A4(n11756), .Y(
        n11752) );
  AND4X1_RVT U11664 ( .A1(n11757), .A2(n11758), .A3(n11350), .A4(n11759), .Y(
        n11756) );
  OR2X1_RVT U11665 ( .A1(n11491), .A2(n11760), .Y(n11350) );
  OR2X1_RVT U11666 ( .A1(n11582), .A2(n136), .Y(n11760) );
  OR2X1_RVT U11667 ( .A1(n11354), .A2(n11761), .Y(n11758) );
  OR2X1_RVT U11668 ( .A1(n12827), .A2(n12830), .Y(n11761) );
  OR2X1_RVT U11669 ( .A1(n11617), .A2(n11762), .Y(n11757) );
  OR2X1_RVT U11670 ( .A1(n11763), .A2(n11391), .Y(n11762) );
  AND2X1_RVT U11671 ( .A1(n12172), .A2(n11491), .Y(n11763) );
  OR2X1_RVT U11672 ( .A1(n11764), .A2(n12178), .Y(n11755) );
  AND2X1_RVT U11673 ( .A1(n11632), .A2(n11704), .Y(n11764) );
  OR2X1_RVT U11674 ( .A1(n136), .A2(n11765), .Y(n11704) );
  OR2X1_RVT U11675 ( .A1(n12151), .A2(n12826), .Y(n11765) );
  OR2X1_RVT U11676 ( .A1(n11421), .A2(n11766), .Y(n11632) );
  OR2X1_RVT U11677 ( .A1(n12824), .A2(n11413), .Y(n11766) );
  OR2X1_RVT U11678 ( .A1(n11767), .A2(n11371), .Y(n11754) );
  AND2X1_RVT U11679 ( .A1(n11768), .A2(n11576), .Y(n11767) );
  OR2X1_RVT U11680 ( .A1(n11477), .A2(n11471), .Y(n11753) );
  AND4X1_RVT U11681 ( .A1(n11769), .A2(n11770), .A3(n11771), .A4(n11772), .Y(
        n11751) );
  AND2X1_RVT U11682 ( .A1(n11773), .A2(n11774), .Y(n11772) );
  OR2X1_RVT U11683 ( .A1(n11775), .A2(n12172), .Y(n11774) );
  AND2X1_RVT U11684 ( .A1(n11776), .A2(n11444), .Y(n11775) );
  AND2X1_RVT U11685 ( .A1(n11777), .A2(n11778), .Y(n11773) );
  OR2X1_RVT U11686 ( .A1(n11779), .A2(n11427), .Y(n11778) );
  AND2X1_RVT U11687 ( .A1(n11398), .A2(n11370), .Y(n11779) );
  OR2X1_RVT U11688 ( .A1(n12832), .A2(n11469), .Y(n11398) );
  OR2X1_RVT U11689 ( .A1(n11780), .A2(n11480), .Y(n11777) );
  AND2X1_RVT U11690 ( .A1(n11672), .A2(n11781), .Y(n11780) );
  OR2X1_RVT U11691 ( .A1(n12833), .A2(n11508), .Y(n11672) );
  OR2X1_RVT U11692 ( .A1(n11782), .A2(n12824), .Y(n11771) );
  AND2X1_RVT U11693 ( .A1(n11375), .A2(n11783), .Y(n11782) );
  OR2X1_RVT U11694 ( .A1(n11511), .A2(n11435), .Y(n11783) );
  OR2X1_RVT U11695 ( .A1(n11414), .A2(n11617), .Y(n11375) );
  OR2X1_RVT U11696 ( .A1(n11784), .A2(n134), .Y(n11770) );
  AND2X1_RVT U11697 ( .A1(n11425), .A2(n11785), .Y(n11784) );
  OR2X1_RVT U11698 ( .A1(n11786), .A2(n12156), .Y(n11785) );
  AND2X1_RVT U11699 ( .A1(n11787), .A2(n11788), .Y(n11786) );
  OR2X1_RVT U11700 ( .A1(n12825), .A2(n11408), .Y(n11788) );
  OR2X1_RVT U11701 ( .A1(n12183), .A2(n11511), .Y(n11425) );
  OR2X1_RVT U11702 ( .A1(n11789), .A2(n11495), .Y(n11769) );
  AND2X1_RVT U11703 ( .A1(n11428), .A2(n11473), .Y(n11789) );
  OR2X1_RVT U11704 ( .A1(n12821), .A2(n11356), .Y(n11473) );
  AND4X1_RVT U11705 ( .A1(n11790), .A2(n11791), .A3(n11792), .A4(n11793), .Y(
        n11750) );
  AND4X1_RVT U11706 ( .A1(n11794), .A2(n11795), .A3(n11796), .A4(n11797), .Y(
        n11793) );
  OR2X1_RVT U11707 ( .A1(n11798), .A2(n12832), .Y(n11797) );
  AND2X1_RVT U11708 ( .A1(n11531), .A2(n11799), .Y(n11798) );
  OR2X1_RVT U11709 ( .A1(n12180), .A2(n11380), .Y(n11799) );
  OR2X1_RVT U11710 ( .A1(n11800), .A2(n11373), .Y(n11796) );
  AND2X1_RVT U11711 ( .A1(n11801), .A2(n11802), .Y(n11800) );
  OR2X1_RVT U11712 ( .A1(n11803), .A2(n11408), .Y(n11802) );
  AND2X1_RVT U11713 ( .A1(n11433), .A2(n11421), .Y(n11803) );
  AND2X1_RVT U11714 ( .A1(n11435), .A2(n11677), .Y(n11801) );
  OR2X1_RVT U11715 ( .A1(n12181), .A2(n11573), .Y(n11677) );
  OR2X1_RVT U11716 ( .A1(n11804), .A2(n12170), .Y(n11795) );
  AND2X1_RVT U11717 ( .A1(n11805), .A2(n11806), .Y(n11804) );
  OR2X1_RVT U11718 ( .A1(n11421), .A2(n11807), .Y(n11806) );
  AND2X1_RVT U11719 ( .A1(n11503), .A2(n11697), .Y(n11805) );
  OR2X1_RVT U11720 ( .A1(n11413), .A2(n11588), .Y(n11697) );
  OR2X1_RVT U11721 ( .A1(n11386), .A2(n11808), .Y(n11503) );
  OR2X1_RVT U11722 ( .A1(n11809), .A2(n11356), .Y(n11794) );
  AND4X1_RVT U11723 ( .A1(n11810), .A2(n11811), .A3(n11812), .A4(n11745), .Y(
        n11809) );
  OR2X1_RVT U11724 ( .A1(n11449), .A2(n11813), .Y(n11745) );
  OR2X1_RVT U11725 ( .A1(n12151), .A2(n11413), .Y(n11813) );
  OR2X1_RVT U11726 ( .A1(n12829), .A2(n11655), .Y(n11811) );
  OR2X1_RVT U11727 ( .A1(n11414), .A2(n11511), .Y(n11810) );
  OR2X1_RVT U11728 ( .A1(n11582), .A2(n11624), .Y(n11792) );
  OR2X1_RVT U11729 ( .A1(n11814), .A2(n12154), .Y(n11791) );
  AND4X1_RVT U11730 ( .A1(n11815), .A2(n11816), .A3(n11458), .A4(n11556), .Y(
        n11814) );
  OR2X1_RVT U11731 ( .A1(n11380), .A2(n11545), .Y(n11556) );
  OR2X1_RVT U11732 ( .A1(n12829), .A2(n134), .Y(n11545) );
  OR2X1_RVT U11733 ( .A1(n11373), .A2(n11437), .Y(n11458) );
  OR2X1_RVT U11734 ( .A1(n12821), .A2(n11808), .Y(n11790) );
  AND4X1_RVT U11735 ( .A1(n11817), .A2(n11818), .A3(n11819), .A4(n11820), .Y(
        n11749) );
  OR2X1_RVT U11736 ( .A1(n12159), .A2(n11821), .Y(n11820) );
  AND2X1_RVT U11737 ( .A1(n11822), .A2(n11823), .Y(n11819) );
  OR2X1_RVT U11738 ( .A1(n12180), .A2(n11576), .Y(n11823) );
  OR2X1_RVT U11739 ( .A1(n11363), .A2(n11437), .Y(n11822) );
  OR2X1_RVT U11740 ( .A1(n136), .A2(n11394), .Y(n11437) );
  OR2X1_RVT U11741 ( .A1(n12183), .A2(n11555), .Y(n11818) );
  OR2X1_RVT U11742 ( .A1(n11430), .A2(n11824), .Y(n11555) );
  AND2X1_RVT U11743 ( .A1(n11825), .A2(n11826), .Y(n11817) );
  OR2X1_RVT U11744 ( .A1(n12152), .A2(n11827), .Y(n11826) );
  OR2X1_RVT U11745 ( .A1(n11433), .A2(n11382), .Y(n11825) );
  OR2X1_RVT U11746 ( .A1(n11356), .A2(n11641), .Y(n11382) );
  AND4X1_RVT U11747 ( .A1(n11829), .A2(n11830), .A3(n11831), .A4(n11832), .Y(
        n11828) );
  AND4X1_RVT U11748 ( .A1(n11833), .A2(n11834), .A3(n11835), .A4(n11836), .Y(
        n11832) );
  AND4X1_RVT U11749 ( .A1(n11569), .A2(n11759), .A3(n11837), .A4(n11838), .Y(
        n11836) );
  OR2X1_RVT U11750 ( .A1(n11839), .A2(n11840), .Y(n11759) );
  OR2X1_RVT U11751 ( .A1(n11354), .A2(n11624), .Y(n11569) );
  OR2X1_RVT U11752 ( .A1(n12830), .A2(n12168), .Y(n11624) );
  AND4X1_RVT U11753 ( .A1(n11827), .A2(n11693), .A3(n11816), .A4(n11351), .Y(
        n11835) );
  OR2X1_RVT U11754 ( .A1(n11841), .A2(n11541), .Y(n11351) );
  OR2X1_RVT U11755 ( .A1(n11356), .A2(n11842), .Y(n11816) );
  OR2X1_RVT U11756 ( .A1(n11389), .A2(n134), .Y(n11693) );
  OR2X1_RVT U11757 ( .A1(n11380), .A2(n11843), .Y(n11827) );
  OR2X1_RVT U11758 ( .A1(n12158), .A2(n12178), .Y(n11843) );
  AND4X1_RVT U11759 ( .A1(n11844), .A2(n11845), .A3(n11846), .A4(n11847), .Y(
        n11834) );
  OR2X1_RVT U11760 ( .A1(n11633), .A2(n11848), .Y(n11847) );
  OR2X1_RVT U11761 ( .A1(n12178), .A2(n11413), .Y(n11848) );
  OR2X1_RVT U11762 ( .A1(n11542), .A2(n11849), .Y(n11846) );
  OR2X1_RVT U11763 ( .A1(n12831), .A2(n11430), .Y(n11849) );
  OR2X1_RVT U11764 ( .A1(n11768), .A2(n11850), .Y(n11845) );
  OR2X1_RVT U11765 ( .A1(n11851), .A2(n11427), .Y(n11850) );
  OR2X1_RVT U11766 ( .A1(n12175), .A2(n11852), .Y(n11844) );
  OR2X1_RVT U11767 ( .A1(n11853), .A2(n12158), .Y(n11852) );
  AND2X1_RVT U11768 ( .A1(n11641), .A2(n11854), .Y(n11853) );
  AND2X1_RVT U11769 ( .A1(n11855), .A2(n11856), .Y(n11833) );
  OR2X1_RVT U11770 ( .A1(n11857), .A2(n11408), .Y(n11856) );
  AND2X1_RVT U11771 ( .A1(n11858), .A2(n11859), .Y(n11857) );
  OR2X1_RVT U11772 ( .A1(n12157), .A2(n11601), .Y(n11859) );
  OR2X1_RVT U11773 ( .A1(n12161), .A2(n11676), .Y(n11858) );
  AND2X1_RVT U11774 ( .A1(n11860), .A2(n11861), .Y(n11855) );
  OR2X1_RVT U11775 ( .A1(n11862), .A2(n11447), .Y(n11861) );
  AND2X1_RVT U11776 ( .A1(n11863), .A2(n11864), .Y(n11862) );
  OR2X1_RVT U11777 ( .A1(n12164), .A2(n144), .Y(n11864) );
  NAND2X1_RVT U11778 ( .A1(n11430), .A2(n12823), .Y(n11863) );
  OR2X1_RVT U11779 ( .A1(n11865), .A2(n136), .Y(n11860) );
  AND2X1_RVT U11780 ( .A1(n11654), .A2(n11531), .Y(n11865) );
  OR2X1_RVT U11781 ( .A1(n11380), .A2(n11866), .Y(n11531) );
  OR2X1_RVT U11782 ( .A1(n12834), .A2(n12153), .Y(n11866) );
  AND4X1_RVT U11783 ( .A1(n11548), .A2(n11867), .A3(n11740), .A4(n11868), .Y(
        n11831) );
  AND4X1_RVT U11784 ( .A1(n11869), .A2(n11870), .A3(n11871), .A4(n11872), .Y(
        n11868) );
  OR2X1_RVT U11785 ( .A1(n11511), .A2(n11432), .Y(n11872) );
  OR2X1_RVT U11786 ( .A1(n11449), .A2(n11478), .Y(n11871) );
  OR2X1_RVT U11787 ( .A1(n12822), .A2(n11703), .Y(n11870) );
  OR2X1_RVT U11788 ( .A1(n11427), .A2(n11409), .Y(n11703) );
  OR2X1_RVT U11789 ( .A1(n12830), .A2(n11491), .Y(n11409) );
  OR2X1_RVT U11790 ( .A1(n12167), .A2(n11532), .Y(n11869) );
  OR2X1_RVT U11791 ( .A1(n11413), .A2(n11641), .Y(n11532) );
  OR2X1_RVT U11792 ( .A1(n12151), .A2(n11617), .Y(n11641) );
  AND2X1_RVT U11793 ( .A1(n11873), .A2(n11874), .Y(n11740) );
  OR2X1_RVT U11794 ( .A1(n11875), .A2(n11480), .Y(n11874) );
  OR2X1_RVT U11795 ( .A1(n12177), .A2(n136), .Y(n11875) );
  OR2X1_RVT U11796 ( .A1(n11876), .A2(n11363), .Y(n11873) );
  OR2X1_RVT U11797 ( .A1(n12821), .A2(n11480), .Y(n11363) );
  OR2X1_RVT U11798 ( .A1(n11377), .A2(n11427), .Y(n11876) );
  OR2X1_RVT U11799 ( .A1(n12159), .A2(n11746), .Y(n11867) );
  AND2X1_RVT U11800 ( .A1(n11877), .A2(n11878), .Y(n11548) );
  OR2X1_RVT U11801 ( .A1(n11431), .A2(n11469), .Y(n11878) );
  OR2X1_RVT U11802 ( .A1(n11879), .A2(n11880), .Y(n11877) );
  AND4X1_RVT U11803 ( .A1(n11881), .A2(n11882), .A3(n11883), .A4(n11884), .Y(
        n11830) );
  OR2X1_RVT U11804 ( .A1(n11885), .A2(n11617), .Y(n11884) );
  AND2X1_RVT U11805 ( .A1(n11886), .A2(n11626), .Y(n11885) );
  OR2X1_RVT U11806 ( .A1(n12165), .A2(n11842), .Y(n11626) );
  OR2X1_RVT U11807 ( .A1(n11887), .A2(n12827), .Y(n11883) );
  AND2X1_RVT U11808 ( .A1(n11554), .A2(n11519), .Y(n11887) );
  OR2X1_RVT U11809 ( .A1(n12821), .A2(n11495), .Y(n11519) );
  OR2X1_RVT U11810 ( .A1(n11888), .A2(n11574), .Y(n11882) );
  AND2X1_RVT U11811 ( .A1(n11889), .A2(n11890), .Y(n11888) );
  OR2X1_RVT U11812 ( .A1(n12154), .A2(n11433), .Y(n11890) );
  AND2X1_RVT U11813 ( .A1(n11891), .A2(n11471), .Y(n11889) );
  OR2X1_RVT U11814 ( .A1(n134), .A2(n11430), .Y(n11891) );
  OR2X1_RVT U11815 ( .A1(n11892), .A2(n11371), .Y(n11881) );
  AND2X1_RVT U11816 ( .A1(n11893), .A2(n11894), .Y(n11892) );
  NAND2X1_RVT U11817 ( .A1(n11356), .A2(n11734), .Y(n11894) );
  AND2X1_RVT U11818 ( .A1(n11895), .A2(n11584), .Y(n11893) );
  OR2X1_RVT U11819 ( .A1(n11517), .A2(n11842), .Y(n11584) );
  OR2X1_RVT U11820 ( .A1(n12174), .A2(n11896), .Y(n11895) );
  AND4X1_RVT U11821 ( .A1(n11897), .A2(n11898), .A3(n11899), .A4(n11900), .Y(
        n11829) );
  OR2X1_RVT U11822 ( .A1(n11901), .A2(n11394), .Y(n11900) );
  AND2X1_RVT U11823 ( .A1(n11902), .A2(n11535), .Y(n11901) );
  AND2X1_RVT U11824 ( .A1(n11903), .A2(n11557), .Y(n11902) );
  OR2X1_RVT U11825 ( .A1(n136), .A2(n11880), .Y(n11557) );
  OR2X1_RVT U11826 ( .A1(n12153), .A2(n11491), .Y(n11880) );
  OR2X1_RVT U11827 ( .A1(n11904), .A2(n12170), .Y(n11899) );
  AND2X1_RVT U11828 ( .A1(n11905), .A2(n11906), .Y(n11904) );
  OR2X1_RVT U11829 ( .A1(n11907), .A2(n12819), .Y(n11906) );
  AND2X1_RVT U11830 ( .A1(n11908), .A2(n11909), .Y(n11907) );
  OR2X1_RVT U11831 ( .A1(n12152), .A2(n11768), .Y(n11909) );
  OR2X1_RVT U11832 ( .A1(n12826), .A2(n11414), .Y(n11908) );
  AND2X1_RVT U11833 ( .A1(n11910), .A2(n11911), .Y(n11905) );
  OR2X1_RVT U11834 ( .A1(n11380), .A2(n11912), .Y(n11910) );
  OR2X1_RVT U11835 ( .A1(n11913), .A2(n11414), .Y(n11898) );
  AND4X1_RVT U11836 ( .A1(n11914), .A2(n11915), .A3(n11916), .A4(n11380), .Y(
        n11913) );
  OR2X1_RVT U11837 ( .A1(n12827), .A2(n11430), .Y(n11916) );
  OR2X1_RVT U11838 ( .A1(n12164), .A2(n11449), .Y(n11915) );
  OR2X1_RVT U11839 ( .A1(n11502), .A2(n11480), .Y(n11914) );
  OR2X1_RVT U11840 ( .A1(n11917), .A2(n11356), .Y(n11897) );
  AND4X1_RVT U11841 ( .A1(n11781), .A2(n11918), .A3(n11579), .A4(n11495), .Y(
        n11917) );
  OR2X1_RVT U11842 ( .A1(n11449), .A2(n11912), .Y(n11579) );
  OR2X1_RVT U11843 ( .A1(n11617), .A2(n11824), .Y(n11918) );
  OR2X1_RVT U11844 ( .A1(n12158), .A2(n11582), .Y(n11781) );
  AND4X1_RVT U11845 ( .A1(n11920), .A2(n11921), .A3(n11922), .A4(n11923), .Y(
        n11919) );
  AND4X1_RVT U11846 ( .A1(n11432), .A2(n11668), .A3(n11924), .A4(n11925), .Y(
        n11923) );
  AND4X1_RVT U11847 ( .A1(n11747), .A2(n11692), .A3(n11837), .A4(n11838), .Y(
        n11925) );
  OR2X1_RVT U11848 ( .A1(n11840), .A2(n11353), .Y(n11838) );
  OR2X1_RVT U11849 ( .A1(n12825), .A2(n11471), .Y(n11353) );
  OR2X1_RVT U11850 ( .A1(n11370), .A2(n11879), .Y(n11837) );
  OR2X1_RVT U11851 ( .A1(n12830), .A2(n12172), .Y(n11879) );
  OR2X1_RVT U11852 ( .A1(n12819), .A2(n11491), .Y(n11370) );
  OR2X1_RVT U11853 ( .A1(n12831), .A2(n11389), .Y(n11692) );
  OR2X1_RVT U11854 ( .A1(n12181), .A2(n12165), .Y(n11389) );
  OR2X1_RVT U11855 ( .A1(n11511), .A2(n11926), .Y(n11747) );
  OR2X1_RVT U11856 ( .A1(n12172), .A2(n11415), .Y(n11926) );
  OR2X1_RVT U11857 ( .A1(n11413), .A2(n11927), .Y(n11924) );
  OR2X1_RVT U11858 ( .A1(n11541), .A2(n12163), .Y(n11927) );
  OR2X1_RVT U11859 ( .A1(n11480), .A2(n11928), .Y(n11668) );
  OR2X1_RVT U11860 ( .A1(n11414), .A2(n12170), .Y(n11928) );
  OR2X1_RVT U11861 ( .A1(n12823), .A2(n11839), .Y(n11432) );
  OR2X1_RVT U11862 ( .A1(n12165), .A2(n11431), .Y(n11839) );
  AND4X1_RVT U11863 ( .A1(n11929), .A2(n11930), .A3(n11931), .A4(n11932), .Y(
        n11922) );
  AND4X1_RVT U11864 ( .A1(n11933), .A2(n11934), .A3(n11935), .A4(n11936), .Y(
        n11932) );
  OR2X1_RVT U11865 ( .A1(n11447), .A2(n11937), .Y(n11936) );
  OR2X1_RVT U11866 ( .A1(n12154), .A2(n11517), .Y(n11937) );
  OR2X1_RVT U11867 ( .A1(n11430), .A2(n11938), .Y(n11935) );
  OR2X1_RVT U11868 ( .A1(n11939), .A2(n11394), .Y(n11938) );
  AND2X1_RVT U11869 ( .A1(n11373), .A2(n11433), .Y(n11939) );
  OR2X1_RVT U11870 ( .A1(n11940), .A2(n11941), .Y(n11934) );
  AND2X1_RVT U11871 ( .A1(n11588), .A2(n11544), .Y(n11940) );
  OR2X1_RVT U11872 ( .A1(n12824), .A2(n144), .Y(n11544) );
  OR2X1_RVT U11873 ( .A1(n12820), .A2(n12175), .Y(n11588) );
  OR2X1_RVT U11874 ( .A1(n11942), .A2(n11428), .Y(n11933) );
  AND2X1_RVT U11875 ( .A1(n11824), .A2(n11943), .Y(n11942) );
  OR2X1_RVT U11876 ( .A1(n12822), .A2(n136), .Y(n11943) );
  OR2X1_RVT U11877 ( .A1(n11944), .A2(n12177), .Y(n11931) );
  AND2X1_RVT U11878 ( .A1(n11815), .A2(n11945), .Y(n11944) );
  OR2X1_RVT U11879 ( .A1(n11421), .A2(n11768), .Y(n11945) );
  OR2X1_RVT U11880 ( .A1(n12158), .A2(n11633), .Y(n11815) );
  OR2X1_RVT U11881 ( .A1(n12826), .A2(n11421), .Y(n11633) );
  OR2X1_RVT U11882 ( .A1(n11946), .A2(n11582), .Y(n11930) );
  AND2X1_RVT U11883 ( .A1(n11535), .A2(n11807), .Y(n11946) );
  OR2X1_RVT U11884 ( .A1(n11391), .A2(n11480), .Y(n11535) );
  OR2X1_RVT U11885 ( .A1(n11947), .A2(n11471), .Y(n11929) );
  AND2X1_RVT U11886 ( .A1(n11434), .A2(n11436), .Y(n11947) );
  AND4X1_RVT U11887 ( .A1(n11948), .A2(n11949), .A3(n11950), .A4(n11951), .Y(
        n11921) );
  AND4X1_RVT U11888 ( .A1(n11952), .A2(n11953), .A3(n11954), .A4(n11955), .Y(
        n11951) );
  OR2X1_RVT U11889 ( .A1(n11956), .A2(n12161), .Y(n11955) );
  AND2X1_RVT U11890 ( .A1(n11362), .A2(n11654), .Y(n11956) );
  OR2X1_RVT U11891 ( .A1(n11511), .A2(n11542), .Y(n11654) );
  OR2X1_RVT U11892 ( .A1(n12164), .A2(n11394), .Y(n11542) );
  OR2X1_RVT U11893 ( .A1(n12168), .A2(n11957), .Y(n11362) );
  OR2X1_RVT U11894 ( .A1(n12151), .A2(n12157), .Y(n11957) );
  OR2X1_RVT U11895 ( .A1(n11958), .A2(n12175), .Y(n11954) );
  AND2X1_RVT U11896 ( .A1(n11671), .A2(n11959), .Y(n11958) );
  OR2X1_RVT U11897 ( .A1(n12180), .A2(n134), .Y(n11959) );
  OR2X1_RVT U11898 ( .A1(n12178), .A2(n11478), .Y(n11671) );
  OR2X1_RVT U11899 ( .A1(n11960), .A2(n12156), .Y(n11953) );
  AND2X1_RVT U11900 ( .A1(n11689), .A2(n11961), .Y(n11960) );
  OR2X1_RVT U11901 ( .A1(n12181), .A2(n11414), .Y(n11961) );
  OR2X1_RVT U11902 ( .A1(n11356), .A2(n11962), .Y(n11689) );
  OR2X1_RVT U11903 ( .A1(n11963), .A2(n11415), .Y(n11952) );
  AND2X1_RVT U11904 ( .A1(n11964), .A2(n11965), .Y(n11963) );
  OR2X1_RVT U11905 ( .A1(n11471), .A2(n12178), .Y(n11965) );
  AND2X1_RVT U11906 ( .A1(n11966), .A2(n11447), .Y(n11964) );
  OR2X1_RVT U11907 ( .A1(n11433), .A2(n11394), .Y(n11447) );
  OR2X1_RVT U11908 ( .A1(n12153), .A2(n11478), .Y(n11966) );
  OR2X1_RVT U11909 ( .A1(n12834), .A2(n11433), .Y(n11478) );
  OR2X1_RVT U11910 ( .A1(n11967), .A2(n11491), .Y(n11950) );
  AND4X1_RVT U11911 ( .A1(n11968), .A2(n11969), .A3(n11644), .A4(n11554), .Y(
        n11967) );
  OR2X1_RVT U11912 ( .A1(n11617), .A2(n11717), .Y(n11554) );
  OR2X1_RVT U11913 ( .A1(n11449), .A2(n11896), .Y(n11644) );
  OR2X1_RVT U11914 ( .A1(n12159), .A2(n12152), .Y(n11896) );
  OR2X1_RVT U11915 ( .A1(n136), .A2(n11371), .Y(n11969) );
  OR2X1_RVT U11916 ( .A1(n134), .A2(n12178), .Y(n11968) );
  OR2X1_RVT U11917 ( .A1(n11970), .A2(n11427), .Y(n11949) );
  AND2X1_RVT U11918 ( .A1(n11971), .A2(n11448), .Y(n11970) );
  AND2X1_RVT U11919 ( .A1(n11903), .A2(n11698), .Y(n11971) );
  OR2X1_RVT U11920 ( .A1(n11972), .A2(n12831), .Y(n11698) );
  AND2X1_RVT U11921 ( .A1(n11469), .A2(n11973), .Y(n11972) );
  OR2X1_RVT U11922 ( .A1(n12156), .A2(n11356), .Y(n11973) );
  OR2X1_RVT U11923 ( .A1(n11517), .A2(n11655), .Y(n11903) );
  OR2X1_RVT U11924 ( .A1(n11502), .A2(n11391), .Y(n11655) );
  OR2X1_RVT U11925 ( .A1(n11974), .A2(n11495), .Y(n11948) );
  AND2X1_RVT U11926 ( .A1(n11975), .A2(n12164), .Y(n11974) );
  AND2X1_RVT U11927 ( .A1(n11976), .A2(n11676), .Y(n11975) );
  OR2X1_RVT U11928 ( .A1(n11517), .A2(n11617), .Y(n11976) );
  AND4X1_RVT U11929 ( .A1(n11977), .A2(n11978), .A3(n11979), .A4(n11980), .Y(
        n11920) );
  AND2X1_RVT U11930 ( .A1(n11981), .A2(n11982), .Y(n11980) );
  OR2X1_RVT U11931 ( .A1(n12827), .A2(n11597), .Y(n11982) );
  OR2X1_RVT U11932 ( .A1(n12172), .A2(n11983), .Y(n11597) );
  OR2X1_RVT U11933 ( .A1(n11413), .A2(n11502), .Y(n11983) );
  AND2X1_RVT U11934 ( .A1(n11984), .A2(n11985), .Y(n11981) );
  OR2X1_RVT U11935 ( .A1(n11386), .A2(n11397), .Y(n11985) );
  OR2X1_RVT U11936 ( .A1(n11430), .A2(n11625), .Y(n11397) );
  OR2X1_RVT U11937 ( .A1(n12823), .A2(n11391), .Y(n11625) );
  OR2X1_RVT U11938 ( .A1(n11433), .A2(n11510), .Y(n11984) );
  OR2X1_RVT U11939 ( .A1(n11421), .A2(n11986), .Y(n11510) );
  OR2X1_RVT U11940 ( .A1(n11421), .A2(n11601), .Y(n11979) );
  OR2X1_RVT U11941 ( .A1(n136), .A2(n12174), .Y(n11601) );
  OR2X1_RVT U11942 ( .A1(n11987), .A2(n11377), .Y(n11978) );
  AND4X1_RVT U11943 ( .A1(n11988), .A2(n11989), .A3(n11990), .A4(n11991), .Y(
        n11987) );
  OR2X1_RVT U11944 ( .A1(n12821), .A2(n11992), .Y(n11990) );
  OR2X1_RVT U11945 ( .A1(n11993), .A2(n12828), .Y(n11992) );
  AND2X1_RVT U11946 ( .A1(n11428), .A2(n11994), .Y(n11993) );
  OR2X1_RVT U11947 ( .A1(n12167), .A2(n11995), .Y(n11989) );
  OR2X1_RVT U11948 ( .A1(n11734), .A2(n11371), .Y(n11995) );
  OR2X1_RVT U11949 ( .A1(n11354), .A2(n11380), .Y(n11988) );
  OR2X1_RVT U11950 ( .A1(n12825), .A2(n11480), .Y(n11380) );
  OR2X1_RVT U11951 ( .A1(n11854), .A2(n11768), .Y(n11977) );
  OR2X1_RVT U11952 ( .A1(n12183), .A2(n11391), .Y(n11768) );
  AND4X1_RVT U11953 ( .A1(n11997), .A2(n11998), .A3(n11999), .A4(n12000), .Y(
        n11996) );
  AND4X1_RVT U11954 ( .A1(n12001), .A2(n12002), .A3(n12003), .A4(n12004), .Y(
        n12000) );
  AND2X1_RVT U11955 ( .A1(n12005), .A2(n12006), .Y(n12004) );
  AND4X1_RVT U11956 ( .A1(n8923), .A2(n8112), .A3(n11016), .A4(n11017), .Y(
        n12006) );
  OR2X1_RVT U11957 ( .A1(n6197), .A2(n10042), .Y(n11017) );
  OR2X1_RVT U11958 ( .A1(n85), .A2(n78), .Y(n10042) );
  OR2X1_RVT U11959 ( .A1(n7030), .A2(n12007), .Y(n11016) );
  OR2X1_RVT U11960 ( .A1(n12876), .A2(n12198), .Y(n12007) );
  OR2X1_RVT U11961 ( .A1(n12149), .A2(n1300), .Y(n7030) );
  OR2X1_RVT U11962 ( .A1(n12926), .A2(n8925), .Y(n8112) );
  OR2X1_RVT U11963 ( .A1(n1312), .A2(n12212), .Y(n8925) );
  OR2X1_RVT U11964 ( .A1(n1332), .A2(n12008), .Y(n8923) );
  OR2X1_RVT U11965 ( .A1(n12211), .A2(n12926), .Y(n12008) );
  AND4X1_RVT U11966 ( .A1(n12009), .A2(n12010), .A3(n12011), .A4(n12012), .Y(
        n12005) );
  OR2X1_RVT U11967 ( .A1(n8061), .A2(n12013), .Y(n12012) );
  OR2X1_RVT U11968 ( .A1(n12014), .A2(n12926), .Y(n12013) );
  OR2X1_RVT U11969 ( .A1(n71), .A2(n8919), .Y(n8061) );
  OR2X1_RVT U11970 ( .A1(n6145), .A2(n12015), .Y(n12011) );
  OR2X1_RVT U11971 ( .A1(n12016), .A2(n12877), .Y(n12015) );
  AND2X1_RVT U11972 ( .A1(n12189), .A2(n8924), .Y(n12016) );
  OR2X1_RVT U11973 ( .A1(n71), .A2(n12868), .Y(n8924) );
  OR2X1_RVT U11974 ( .A1(n12017), .A2(n8056), .Y(n12010) );
  OR2X1_RVT U11975 ( .A1(n8919), .A2(n12212), .Y(n8056) );
  AND2X1_RVT U11976 ( .A1(n8122), .A2(n12018), .Y(n12017) );
  OR2X1_RVT U11977 ( .A1(n1328), .A2(n12191), .Y(n12018) );
  OR2X1_RVT U11978 ( .A1(n12019), .A2(n6128), .Y(n12009) );
  AND2X1_RVT U11979 ( .A1(n8946), .A2(n8088), .Y(n12019) );
  OR2X1_RVT U11980 ( .A1(n1312), .A2(n1300), .Y(n8946) );
  AND4X1_RVT U11981 ( .A1(n12020), .A2(n12021), .A3(n12022), .A4(n12023), .Y(
        n12003) );
  OR2X1_RVT U11982 ( .A1(n12024), .A2(n1332), .Y(n12023) );
  AND2X1_RVT U11983 ( .A1(n1342), .A2(n12025), .Y(n12024) );
  OR2X1_RVT U11984 ( .A1(n6172), .A2(n12026), .Y(n12025) );
  OR2X1_RVT U11985 ( .A1(n1361), .A2(n12871), .Y(n12026) );
  OR2X1_RVT U11986 ( .A1(n1350), .A2(n1334), .Y(n6172) );
  OR2X1_RVT U11987 ( .A1(n12211), .A2(n1388), .Y(n1342) );
  OR2X1_RVT U11988 ( .A1(n12027), .A2(n8919), .Y(n12022) );
  OR2X1_RVT U11989 ( .A1(n12873), .A2(n1312), .Y(n8919) );
  AND2X1_RVT U11990 ( .A1(n6138), .A2(n7032), .Y(n12027) );
  OR2X1_RVT U11991 ( .A1(n71), .A2(n1331), .Y(n7032) );
  OR2X1_RVT U11992 ( .A1(n12928), .A2(n10084), .Y(n6138) );
  OR2X1_RVT U11993 ( .A1(n12028), .A2(n76), .Y(n12021) );
  AND2X1_RVT U11994 ( .A1(n1304), .A2(n10061), .Y(n12028) );
  OR2X1_RVT U11995 ( .A1(n85), .A2(n11030), .Y(n10061) );
  OR2X1_RVT U11996 ( .A1(n12874), .A2(n12211), .Y(n11030) );
  OR2X1_RVT U11997 ( .A1(n12192), .A2(n6197), .Y(n1304) );
  OR2X1_RVT U11998 ( .A1(n12029), .A2(n1300), .Y(n12020) );
  AND2X1_RVT U11999 ( .A1(n7049), .A2(n11074), .Y(n12029) );
  OR2X1_RVT U12000 ( .A1(n12206), .A2(n12030), .Y(n11074) );
  OR2X1_RVT U12001 ( .A1(n12928), .A2(n83), .Y(n12030) );
  OR2X1_RVT U12002 ( .A1(n6198), .A2(n12031), .Y(n7049) );
  OR2X1_RVT U12003 ( .A1(n12874), .A2(n12149), .Y(n12031) );
  OR2X1_RVT U12004 ( .A1(n12032), .A2(n12198), .Y(n12002) );
  AND2X1_RVT U12005 ( .A1(n12033), .A2(n12034), .Y(n12032) );
  OR2X1_RVT U12006 ( .A1(n12035), .A2(n12211), .Y(n12034) );
  AND2X1_RVT U12007 ( .A1(n1314), .A2(n72), .Y(n12035) );
  AND2X1_RVT U12008 ( .A1(n6155), .A2(n1323), .Y(n12033) );
  OR2X1_RVT U12009 ( .A1(n12206), .A2(n12036), .Y(n6155) );
  OR2X1_RVT U12010 ( .A1(n7034), .A2(n12185), .Y(n12036) );
  AND2X1_RVT U12011 ( .A1(n12037), .A2(n12038), .Y(n12001) );
  OR2X1_RVT U12012 ( .A1(n12039), .A2(n8063), .Y(n12038) );
  AND2X1_RVT U12013 ( .A1(n12040), .A2(n12041), .Y(n12039) );
  OR2X1_RVT U12014 ( .A1(n6999), .A2(n6192), .Y(n12041) );
  OR2X1_RVT U12015 ( .A1(n12188), .A2(n72), .Y(n6192) );
  XOR2X1_RVT U12016 ( .A1(n12192), .A2(n12149), .Y(n6999) );
  OR2X1_RVT U12017 ( .A1(n12926), .A2(n6989), .Y(n12040) );
  OR2X1_RVT U12018 ( .A1(n12042), .A2(n1350), .Y(n12037) );
  AND2X1_RVT U12019 ( .A1(n1401), .A2(n8082), .Y(n12042) );
  OR2X1_RVT U12020 ( .A1(n78), .A2(n10084), .Y(n8082) );
  OR2X1_RVT U12021 ( .A1(n12212), .A2(n6128), .Y(n1401) );
  OR2X1_RVT U12022 ( .A1(n8063), .A2(n12209), .Y(n6128) );
  OR2X1_RVT U12023 ( .A1(n12872), .A2(n71), .Y(n1356) );
  AND4X1_RVT U12024 ( .A1(n12043), .A2(n12044), .A3(n12045), .A4(n12046), .Y(
        n11999) );
  AND4X1_RVT U12025 ( .A1(n12047), .A2(n12048), .A3(n12049), .A4(n12050), .Y(
        n12046) );
  OR2X1_RVT U12026 ( .A1(n12196), .A2(n6182), .Y(n12050) );
  OR2X1_RVT U12027 ( .A1(n6198), .A2(n12051), .Y(n6182) );
  OR2X1_RVT U12028 ( .A1(n1325), .A2(n1350), .Y(n12051) );
  OR2X1_RVT U12029 ( .A1(n12868), .A2(n6132), .Y(n6198) );
  OR2X1_RVT U12030 ( .A1(n7034), .A2(n10071), .Y(n12049) );
  OR2X1_RVT U12031 ( .A1(n12206), .A2(n11018), .Y(n10071) );
  OR2X1_RVT U12032 ( .A1(n12926), .A2(n12192), .Y(n11018) );
  OR2X1_RVT U12033 ( .A1(n12870), .A2(n8937), .Y(n12048) );
  OR2X1_RVT U12034 ( .A1(n12195), .A2(n8088), .Y(n8937) );
  OR2X1_RVT U12035 ( .A1(n7034), .A2(n12876), .Y(n8088) );
  OR2X1_RVT U12036 ( .A1(n73), .A2(n7044), .Y(n12047) );
  OR2X1_RVT U12037 ( .A1(n12201), .A2(n8917), .Y(n7044) );
  OR2X1_RVT U12038 ( .A1(n12928), .A2(n1341), .Y(n8917) );
  OR2X1_RVT U12039 ( .A1(n1323), .A2(n1391), .Y(n12045) );
  OR2X1_RVT U12040 ( .A1(n6132), .A2(n12192), .Y(n1391) );
  OR2X1_RVT U12041 ( .A1(n12206), .A2(n10095), .Y(n12044) );
  OR2X1_RVT U12042 ( .A1(n12870), .A2(n1385), .Y(n10095) );
  OR2X1_RVT U12043 ( .A1(n71), .A2(n12208), .Y(n1385) );
  OR2X1_RVT U12044 ( .A1(n1307), .A2(n8912), .Y(n12043) );
  OR2X1_RVT U12045 ( .A1(n12877), .A2(n10056), .Y(n8912) );
  OR2X1_RVT U12046 ( .A1(n12928), .A2(n6132), .Y(n10056) );
  OR2X1_RVT U12047 ( .A1(n12184), .A2(n8063), .Y(n6132) );
  AND4X1_RVT U12048 ( .A1(n12052), .A2(n12053), .A3(n12054), .A4(n12055), .Y(
        n11998) );
  OR2X1_RVT U12049 ( .A1(n12056), .A2(n12189), .Y(n12055) );
  AND2X1_RVT U12050 ( .A1(n12057), .A2(n12058), .Y(n12056) );
  OR2X1_RVT U12051 ( .A1(n69), .A2(n8122), .Y(n12058) );
  OR2X1_RVT U12052 ( .A1(n12867), .A2(n76), .Y(n8122) );
  AND2X1_RVT U12053 ( .A1(n1302), .A2(n1323), .Y(n12057) );
  OR2X1_RVT U12054 ( .A1(n1334), .A2(n1365), .Y(n1323) );
  OR2X1_RVT U12055 ( .A1(n6139), .A2(n72), .Y(n1302) );
  AND2X1_RVT U12056 ( .A1(n73), .A2(n12193), .Y(n8901) );
  OR2X1_RVT U12057 ( .A1(n12184), .A2(n12870), .Y(n6139) );
  OR2X1_RVT U12058 ( .A1(n12059), .A2(n12867), .Y(n12054) );
  AND4X1_RVT U12059 ( .A1(n12060), .A2(n10094), .A3(n8887), .A4(n6196), .Y(
        n12059) );
  OR2X1_RVT U12060 ( .A1(n12189), .A2(n1365), .Y(n6196) );
  OR2X1_RVT U12061 ( .A1(n12928), .A2(n1346), .Y(n8887) );
  OR2X1_RVT U12062 ( .A1(n12201), .A2(n1388), .Y(n1346) );
  OR2X1_RVT U12063 ( .A1(n12209), .A2(n7006), .Y(n10094) );
  OR2X1_RVT U12064 ( .A1(n12871), .A2(n69), .Y(n7006) );
  OR2X1_RVT U12065 ( .A1(n12196), .A2(n1375), .Y(n6145) );
  OR2X1_RVT U12066 ( .A1(n78), .A2(n1365), .Y(n12060) );
  OR2X1_RVT U12067 ( .A1(n69), .A2(n1350), .Y(n1365) );
  OR2X1_RVT U12068 ( .A1(n6197), .A2(n6143), .Y(n12053) );
  OR2X1_RVT U12069 ( .A1(n83), .A2(n12185), .Y(n6143) );
  AND2X1_RVT U12070 ( .A1(n12191), .A2(n85), .Y(n12014) );
  OR2X1_RVT U12071 ( .A1(n12872), .A2(n8055), .Y(n6197) );
  OR2X1_RVT U12072 ( .A1(n1331), .A2(n6989), .Y(n12052) );
  OR2X1_RVT U12073 ( .A1(n1300), .A2(n1388), .Y(n6989) );
  OR2X1_RVT U12074 ( .A1(n73), .A2(n12194), .Y(n1388) );
  OR2X1_RVT U12075 ( .A1(n71), .A2(n12188), .Y(n1300) );
  OR2X1_RVT U12076 ( .A1(n12198), .A2(n76), .Y(n1331) );
  AND2X1_RVT U12077 ( .A1(n12186), .A2(n12928), .Y(n1328) );
  AND4X1_RVT U12078 ( .A1(n12061), .A2(n12062), .A3(n12063), .A4(n12064), .Y(
        n11997) );
  OR2X1_RVT U12079 ( .A1(n1370), .A2(n7008), .Y(n12064) );
  OR2X1_RVT U12080 ( .A1(n12194), .A2(n12201), .Y(n7008) );
  OR2X1_RVT U12081 ( .A1(n12187), .A2(n7034), .Y(n1307) );
  OR2X1_RVT U12082 ( .A1(n12869), .A2(n12926), .Y(n1370) );
  OR2X1_RVT U12083 ( .A1(n12150), .A2(n1375), .Y(n1314) );
  OR2X1_RVT U12084 ( .A1(n78), .A2(n8892), .Y(n12063) );
  OR2X1_RVT U12085 ( .A1(n12198), .A2(n12065), .Y(n8892) );
  OR2X1_RVT U12086 ( .A1(n73), .A2(n7034), .Y(n12065) );
  OR2X1_RVT U12087 ( .A1(n12867), .A2(n85), .Y(n1341) );
  AND2X1_RVT U12088 ( .A1(n12185), .A2(n12195), .Y(n8065) );
  OR2X1_RVT U12089 ( .A1(n12150), .A2(n10062), .Y(n12062) );
  OR2X1_RVT U12090 ( .A1(n6200), .A2(n1332), .Y(n10062) );
  OR2X1_RVT U12091 ( .A1(n8063), .A2(n12192), .Y(n1332) );
  OR2X1_RVT U12092 ( .A1(n1325), .A2(n12877), .Y(n6200) );
  AND2X1_RVT U12093 ( .A1(n1312), .A2(n1350), .Y(n7012) );
  OR2X1_RVT U12094 ( .A1(n7034), .A2(n12189), .Y(n1325) );
  XOR2X1_RVT U12095 ( .A1(key[100]), .A2(state[100]), .Y(n1334) );
  OR2X1_RVT U12096 ( .A1(n11041), .A2(n8055), .Y(n12061) );
  OR2X1_RVT U12097 ( .A1(n12873), .A2(n69), .Y(n8055) );
  AND2X1_RVT U12098 ( .A1(n73), .A2(n71), .Y(n1361) );
  XOR2X1_RVT U12099 ( .A1(key[103]), .A2(state[103]), .Y(n7034) );
  XOR2X1_RVT U12100 ( .A1(key[102]), .A2(state[102]), .Y(n1312) );
  XOR2X1_RVT U12101 ( .A1(key[101]), .A2(state[101]), .Y(n1350) );
  OR2X1_RVT U12102 ( .A1(n12186), .A2(n10084), .Y(n11041) );
  OR2X1_RVT U12103 ( .A1(n12188), .A2(n12869), .Y(n10084) );
  AND2X1_RVT U12104 ( .A1(n8063), .A2(n12868), .Y(n8100) );
  XOR2X1_RVT U12105 ( .A1(key[98]), .A2(state[98]), .Y(n6183) );
  XOR2X1_RVT U12106 ( .A1(key[96]), .A2(state[96]), .Y(n8063) );
  XOR2X1_RVT U12107 ( .A1(key[99]), .A2(state[99]), .Y(n1309) );
  XOR2X1_RVT U12108 ( .A1(key[97]), .A2(state[97]), .Y(n1375) );
  AND4X1_RVT U12109 ( .A1(n12067), .A2(n12068), .A3(n12069), .A4(n12070), .Y(
        n12066) );
  AND4X1_RVT U12110 ( .A1(n12071), .A2(n12072), .A3(n12073), .A4(n12074), .Y(
        n12070) );
  AND4X1_RVT U12111 ( .A1(n12075), .A2(n12076), .A3(n12077), .A4(n12078), .Y(
        n12074) );
  OR2X1_RVT U12112 ( .A1(n11842), .A2(n11986), .Y(n12078) );
  OR2X1_RVT U12113 ( .A1(n12824), .A2(n12177), .Y(n11986) );
  OR2X1_RVT U12114 ( .A1(n12151), .A2(n12161), .Y(n11842) );
  OR2X1_RVT U12115 ( .A1(n12079), .A2(n11428), .Y(n12077) );
  AND2X1_RVT U12116 ( .A1(n11374), .A2(n11941), .Y(n12079) );
  OR2X1_RVT U12117 ( .A1(n136), .A2(n12080), .Y(n11374) );
  OR2X1_RVT U12118 ( .A1(n12151), .A2(n12821), .Y(n12080) );
  OR2X1_RVT U12119 ( .A1(n12081), .A2(n11356), .Y(n12076) );
  OR2X1_RVT U12120 ( .A1(n12165), .A2(n11517), .Y(n11356) );
  AND2X1_RVT U12121 ( .A1(n11492), .A2(n12082), .Y(n12081) );
  OR2X1_RVT U12122 ( .A1(n11371), .A2(n11573), .Y(n12082) );
  OR2X1_RVT U12123 ( .A1(n12169), .A2(n12157), .Y(n11371) );
  OR2X1_RVT U12124 ( .A1(n11617), .A2(n12083), .Y(n11492) );
  OR2X1_RVT U12125 ( .A1(n12832), .A2(n12172), .Y(n12083) );
  OR2X1_RVT U12126 ( .A1(n12084), .A2(n11415), .Y(n12075) );
  AND2X1_RVT U12127 ( .A1(n11812), .A2(n12085), .Y(n12084) );
  OR2X1_RVT U12128 ( .A1(n12086), .A2(n12821), .Y(n12085) );
  AND2X1_RVT U12129 ( .A1(n11471), .A2(n11824), .Y(n12086) );
  OR2X1_RVT U12130 ( .A1(n12829), .A2(n11433), .Y(n11824) );
  OR2X1_RVT U12131 ( .A1(n12178), .A2(n12087), .Y(n11812) );
  OR2X1_RVT U12132 ( .A1(n12834), .A2(n12830), .Y(n12087) );
  OR2X1_RVT U12133 ( .A1(n12088), .A2(n12156), .Y(n12073) );
  AND2X1_RVT U12134 ( .A1(n12089), .A2(n12090), .Y(n12088) );
  OR2X1_RVT U12135 ( .A1(n12091), .A2(n11517), .Y(n12090) );
  AND2X1_RVT U12136 ( .A1(n11582), .A2(n12092), .Y(n12091) );
  OR2X1_RVT U12137 ( .A1(n11373), .A2(n11495), .Y(n12089) );
  OR2X1_RVT U12138 ( .A1(n12170), .A2(n11431), .Y(n11495) );
  OR2X1_RVT U12139 ( .A1(n12093), .A2(n12830), .Y(n12072) );
  AND2X1_RVT U12140 ( .A1(n11587), .A2(n11746), .Y(n12093) );
  OR2X1_RVT U12141 ( .A1(n12168), .A2(n12094), .Y(n11746) );
  OR2X1_RVT U12142 ( .A1(n11427), .A2(n12157), .Y(n12094) );
  OR2X1_RVT U12143 ( .A1(n11373), .A2(n11854), .Y(n11587) );
  OR2X1_RVT U12144 ( .A1(n12157), .A2(n12172), .Y(n11854) );
  OR2X1_RVT U12145 ( .A1(n12095), .A2(n12154), .Y(n12071) );
  AND2X1_RVT U12146 ( .A1(n11627), .A2(n12096), .Y(n12095) );
  OR2X1_RVT U12147 ( .A1(n11841), .A2(n11421), .Y(n12096) );
  OR2X1_RVT U12148 ( .A1(n11480), .A2(n11962), .Y(n11627) );
  OR2X1_RVT U12149 ( .A1(n12829), .A2(n136), .Y(n11962) );
  AND2X1_RVT U12150 ( .A1(n12158), .A2(n12832), .Y(n11723) );
  AND4X1_RVT U12151 ( .A1(n12097), .A2(n12098), .A3(n12099), .A4(n12100), .Y(
        n12069) );
  AND4X1_RVT U12152 ( .A1(n12101), .A2(n12102), .A3(n12103), .A4(n12104), .Y(
        n12100) );
  OR2X1_RVT U12153 ( .A1(n12105), .A2(n12163), .Y(n12104) );
  AND2X1_RVT U12154 ( .A1(n11614), .A2(n11685), .Y(n12105) );
  OR2X1_RVT U12155 ( .A1(n11430), .A2(n11941), .Y(n11685) );
  OR2X1_RVT U12156 ( .A1(n12832), .A2(n11427), .Y(n11941) );
  OR2X1_RVT U12157 ( .A1(n12819), .A2(n12153), .Y(n11430) );
  OR2X1_RVT U12158 ( .A1(n12154), .A2(n11717), .Y(n11614) );
  OR2X1_RVT U12159 ( .A1(n12158), .A2(n12172), .Y(n11717) );
  OR2X1_RVT U12160 ( .A1(n12106), .A2(n12828), .Y(n12103) );
  AND2X1_RVT U12161 ( .A1(n11776), .A2(n12107), .Y(n12106) );
  OR2X1_RVT U12162 ( .A1(n11734), .A2(n11444), .Y(n12107) );
  OR2X1_RVT U12163 ( .A1(n11617), .A2(n12108), .Y(n11444) );
  OR2X1_RVT U12164 ( .A1(n12183), .A2(n12159), .Y(n12108) );
  OR2X1_RVT U12165 ( .A1(n12167), .A2(n12109), .Y(n11776) );
  OR2X1_RVT U12166 ( .A1(n11617), .A2(n11413), .Y(n12109) );
  OR2X1_RVT U12167 ( .A1(n12110), .A2(n12834), .Y(n12102) );
  AND2X1_RVT U12168 ( .A1(n11722), .A2(n11651), .Y(n12110) );
  OR2X1_RVT U12169 ( .A1(n11433), .A2(n11469), .Y(n11651) );
  OR2X1_RVT U12170 ( .A1(n12826), .A2(n11617), .Y(n11469) );
  OR2X1_RVT U12171 ( .A1(n11841), .A2(n11449), .Y(n11722) );
  OR2X1_RVT U12172 ( .A1(n12164), .A2(n12831), .Y(n11841) );
  OR2X1_RVT U12173 ( .A1(n12111), .A2(n11491), .Y(n12101) );
  AND2X1_RVT U12174 ( .A1(n12112), .A2(n12113), .Y(n12111) );
  OR2X1_RVT U12175 ( .A1(n11413), .A2(n11840), .Y(n12113) );
  OR2X1_RVT U12176 ( .A1(n12828), .A2(n144), .Y(n11840) );
  AND2X1_RVT U12177 ( .A1(n12114), .A2(n11708), .Y(n12112) );
  OR2X1_RVT U12178 ( .A1(n11421), .A2(n12115), .Y(n11708) );
  OR2X1_RVT U12179 ( .A1(n12180), .A2(n12159), .Y(n12115) );
  OR2X1_RVT U12180 ( .A1(n11477), .A2(n11414), .Y(n12099) );
  OR2X1_RVT U12181 ( .A1(n12821), .A2(n11373), .Y(n11477) );
  OR2X1_RVT U12182 ( .A1(n12116), .A2(n11377), .Y(n12098) );
  AND2X1_RVT U12183 ( .A1(n12117), .A2(n11558), .Y(n12116) );
  AND2X1_RVT U12184 ( .A1(n12118), .A2(n12119), .Y(n11558) );
  OR2X1_RVT U12185 ( .A1(n12168), .A2(n11582), .Y(n12119) );
  OR2X1_RVT U12186 ( .A1(n11480), .A2(n11354), .Y(n12118) );
  OR2X1_RVT U12187 ( .A1(n12153), .A2(n11427), .Y(n11354) );
  AND2X1_RVT U12188 ( .A1(n12120), .A2(n11744), .Y(n12117) );
  OR2X1_RVT U12189 ( .A1(n11511), .A2(n11994), .Y(n11744) );
  OR2X1_RVT U12190 ( .A1(n12823), .A2(n134), .Y(n11994) );
  OR2X1_RVT U12191 ( .A1(n11373), .A2(n11540), .Y(n12120) );
  OR2X1_RVT U12192 ( .A1(n12152), .A2(n12121), .Y(n11540) );
  OR2X1_RVT U12193 ( .A1(n12819), .A2(n12181), .Y(n12121) );
  OR2X1_RVT U12194 ( .A1(n12122), .A2(n12819), .Y(n12097) );
  AND4X1_RVT U12195 ( .A1(n12123), .A2(n12124), .A3(n12125), .A4(n11886), .Y(
        n12122) );
  OR2X1_RVT U12196 ( .A1(n11427), .A2(n11807), .Y(n11886) );
  OR2X1_RVT U12197 ( .A1(n12824), .A2(n12830), .Y(n11807) );
  OR2X1_RVT U12198 ( .A1(n11427), .A2(n12126), .Y(n12125) );
  OR2X1_RVT U12199 ( .A1(n12158), .A2(n12163), .Y(n12126) );
  OR2X1_RVT U12200 ( .A1(n12829), .A2(n11386), .Y(n11427) );
  OR2X1_RVT U12201 ( .A1(n12127), .A2(n11508), .Y(n12124) );
  OR2X1_RVT U12202 ( .A1(n12152), .A2(n11352), .Y(n11508) );
  AND2X1_RVT U12203 ( .A1(n11491), .A2(n12128), .Y(n12127) );
  OR2X1_RVT U12204 ( .A1(n12827), .A2(n11391), .Y(n12128) );
  OR2X1_RVT U12205 ( .A1(n12823), .A2(n12163), .Y(n11491) );
  OR2X1_RVT U12206 ( .A1(n12825), .A2(n12092), .Y(n12123) );
  OR2X1_RVT U12207 ( .A1(n12829), .A2(n11431), .Y(n12092) );
  OR2X1_RVT U12208 ( .A1(n11377), .A2(n134), .Y(n11431) );
  AND4X1_RVT U12209 ( .A1(n12129), .A2(n12130), .A3(n12131), .A4(n12132), .Y(
        n12068) );
  AND4X1_RVT U12210 ( .A1(n12133), .A2(n12134), .A3(n12135), .A4(n12136), .Y(
        n12132) );
  OR2X1_RVT U12211 ( .A1(n11449), .A2(n11576), .Y(n12136) );
  OR2X1_RVT U12212 ( .A1(n12165), .A2(n11471), .Y(n11576) );
  OR2X1_RVT U12213 ( .A1(n12169), .A2(n11617), .Y(n11449) );
  OR2X1_RVT U12214 ( .A1(n11436), .A2(n11912), .Y(n12135) );
  OR2X1_RVT U12215 ( .A1(n12833), .A2(n12152), .Y(n11912) );
  OR2X1_RVT U12216 ( .A1(n11502), .A2(n11428), .Y(n11436) );
  OR2X1_RVT U12217 ( .A1(n11421), .A2(n11448), .Y(n12134) );
  OR2X1_RVT U12218 ( .A1(n12161), .A2(n12174), .Y(n11448) );
  OR2X1_RVT U12219 ( .A1(n12151), .A2(n12820), .Y(n11421) );
  OR2X1_RVT U12220 ( .A1(n144), .A2(n11787), .Y(n12133) );
  OR2X1_RVT U12221 ( .A1(n12159), .A2(n11574), .Y(n11787) );
  OR2X1_RVT U12222 ( .A1(n11391), .A2(n11821), .Y(n12131) );
  OR2X1_RVT U12223 ( .A1(n144), .A2(n12137), .Y(n11821) );
  OR2X1_RVT U12224 ( .A1(n12826), .A2(n12172), .Y(n12137) );
  AND2X1_RVT U12225 ( .A1(n12153), .A2(n12156), .Y(n11851) );
  OR2X1_RVT U12226 ( .A1(n11433), .A2(n11381), .Y(n12130) );
  OR2X1_RVT U12227 ( .A1(n12181), .A2(n12138), .Y(n11381) );
  OR2X1_RVT U12228 ( .A1(n12827), .A2(n12819), .Y(n12138) );
  OR2X1_RVT U12229 ( .A1(n12158), .A2(n11413), .Y(n11433) );
  OR2X1_RVT U12230 ( .A1(n11480), .A2(n12114), .Y(n12129) );
  OR2X1_RVT U12231 ( .A1(n12154), .A2(n11435), .Y(n12114) );
  OR2X1_RVT U12232 ( .A1(n12829), .A2(n12830), .Y(n11435) );
  AND4X1_RVT U12233 ( .A1(n12139), .A2(n11546), .A3(n12140), .A4(n12141), .Y(
        n12067) );
  OR2X1_RVT U12234 ( .A1(n12158), .A2(n11991), .Y(n12141) );
  OR2X1_RVT U12235 ( .A1(n12825), .A2(n11541), .Y(n11991) );
  OR2X1_RVT U12236 ( .A1(n12156), .A2(n11582), .Y(n11541) );
  OR2X1_RVT U12237 ( .A1(n12151), .A2(n11408), .Y(n11582) );
  AND2X1_RVT U12238 ( .A1(n12142), .A2(n12143), .Y(n12140) );
  OR2X1_RVT U12239 ( .A1(n12180), .A2(n11911), .Y(n12143) );
  OR2X1_RVT U12240 ( .A1(n11480), .A2(n11573), .Y(n11911) );
  OR2X1_RVT U12241 ( .A1(n12158), .A2(n12152), .Y(n11573) );
  OR2X1_RVT U12242 ( .A1(n12153), .A2(n11369), .Y(n11408) );
  OR2X1_RVT U12243 ( .A1(n12832), .A2(n11642), .Y(n12142) );
  OR2X1_RVT U12244 ( .A1(n12177), .A2(n11676), .Y(n11642) );
  OR2X1_RVT U12245 ( .A1(n12824), .A2(n12819), .Y(n11676) );
  OR2X1_RVT U12246 ( .A1(n12822), .A2(n12169), .Y(n11352) );
  AND2X1_RVT U12247 ( .A1(n12144), .A2(n12145), .Y(n11546) );
  OR2X1_RVT U12248 ( .A1(n11428), .A2(n11414), .Y(n12145) );
  OR2X1_RVT U12249 ( .A1(n12831), .A2(n11386), .Y(n11414) );
  AND2X1_RVT U12250 ( .A1(n11413), .A2(n11377), .Y(n11466) );
  OR2X1_RVT U12251 ( .A1(n12164), .A2(n11480), .Y(n11428) );
  OR2X1_RVT U12252 ( .A1(n12820), .A2(n11517), .Y(n11480) );
  OR2X1_RVT U12253 ( .A1(n12146), .A2(n11471), .Y(n12144) );
  OR2X1_RVT U12254 ( .A1(n12158), .A2(n134), .Y(n11471) );
  AND2X1_RVT U12255 ( .A1(n12833), .A2(n12151), .Y(n11734) );
  OR2X1_RVT U12256 ( .A1(n12157), .A2(n11574), .Y(n12146) );
  OR2X1_RVT U12257 ( .A1(n12829), .A2(n12174), .Y(n11574) );
  AND2X1_RVT U12258 ( .A1(n12147), .A2(n12148), .Y(n12139) );
  OR2X1_RVT U12259 ( .A1(n11394), .A2(n11727), .Y(n12148) );
  OR2X1_RVT U12260 ( .A1(n12159), .A2(n11434), .Y(n11727) );
  OR2X1_RVT U12261 ( .A1(n12174), .A2(n11511), .Y(n11434) );
  OR2X1_RVT U12262 ( .A1(n12154), .A2(n12157), .Y(n11511) );
  OR2X1_RVT U12263 ( .A1(n12826), .A2(n12824), .Y(n11373) );
  OR2X1_RVT U12264 ( .A1(n12834), .A2(n12828), .Y(n11394) );
  XOR2X1_RVT U12265 ( .A1(key[76]), .A2(state[76]), .Y(n11369) );
  OR2X1_RVT U12266 ( .A1(n11386), .A2(n11515), .Y(n12147) );
  OR2X1_RVT U12267 ( .A1(n11617), .A2(n11808), .Y(n11515) );
  OR2X1_RVT U12268 ( .A1(n12161), .A2(n11415), .Y(n11808) );
  OR2X1_RVT U12269 ( .A1(n12827), .A2(n11517), .Y(n11415) );
  XOR2X1_RVT U12270 ( .A1(key[74]), .A2(state[74]), .Y(n11517) );
  XOR2X1_RVT U12271 ( .A1(key[75]), .A2(state[75]), .Y(n11451) );
  OR2X1_RVT U12272 ( .A1(n12832), .A2(n12159), .Y(n11391) );
  XOR2X1_RVT U12273 ( .A1(key[77]), .A2(state[77]), .Y(n11377) );
  XOR2X1_RVT U12274 ( .A1(key[78]), .A2(state[78]), .Y(n11413) );
  OR2X1_RVT U12275 ( .A1(n12822), .A2(n12157), .Y(n11617) );
  XOR2X1_RVT U12276 ( .A1(key[72]), .A2(state[72]), .Y(n11392) );
  XOR2X1_RVT U12277 ( .A1(key[73]), .A2(state[73]), .Y(n11502) );
  XOR2X1_RVT U12278 ( .A1(key[79]), .A2(state[79]), .Y(n11386) );
  INVX1_RVT U12279 ( .A(n12196), .Y(n12149) );
  INVX1_RVT U12280 ( .A(n12195), .Y(n12150) );
  INVX1_RVT U12281 ( .A(n11386), .Y(n12151) );
  INVX1_RVT U12282 ( .A(n12151), .Y(n12152) );
  XOR2X1_RVT U12283 ( .A1(key[73]), .A2(state[73]), .Y(n12153) );
  XOR2X1_RVT U12284 ( .A1(key[73]), .A2(state[73]), .Y(n12154) );
  INVX1_RVT U12285 ( .A(n11392), .Y(n12155) );
  INVX1_RVT U12286 ( .A(n12155), .Y(n12156) );
  INVX1_RVT U12287 ( .A(n12155), .Y(n12157) );
  INVX1_RVT U12288 ( .A(n11377), .Y(n12158) );
  INVX1_RVT U12289 ( .A(n12158), .Y(n12159) );
  INVX1_RVT U12290 ( .A(n11391), .Y(n12160) );
  INVX1_RVT U12291 ( .A(n12160), .Y(n12161) );
  INVX1_RVT U12292 ( .A(n11451), .Y(n12162) );
  INVX1_RVT U12293 ( .A(n12162), .Y(n12163) );
  INVX1_RVT U12294 ( .A(n12162), .Y(n12164) );
  INVX1_RVT U12295 ( .A(n12162), .Y(n12165) );
  INVX1_RVT U12296 ( .A(n11415), .Y(n12166) );
  INVX1_RVT U12297 ( .A(n12166), .Y(n12167) );
  INVX1_RVT U12298 ( .A(n12166), .Y(n12168) );
  INVX1_RVT U12299 ( .A(n12828), .Y(n12169) );
  INVX1_RVT U12300 ( .A(n12829), .Y(n12170) );
  INVX1_RVT U12301 ( .A(n11394), .Y(n12171) );
  INVX1_RVT U12302 ( .A(n12171), .Y(n12172) );
  INVX1_RVT U12303 ( .A(n11373), .Y(n12173) );
  INVX1_RVT U12304 ( .A(n12173), .Y(n12174) );
  INVX1_RVT U12305 ( .A(n12173), .Y(n12175) );
  INVX1_RVT U12306 ( .A(n11352), .Y(n12176) );
  INVX1_RVT U12307 ( .A(n12176), .Y(n12177) );
  INVX1_RVT U12308 ( .A(n12176), .Y(n12178) );
  INVX1_RVT U12309 ( .A(n11408), .Y(n12179) );
  INVX1_RVT U12310 ( .A(n12179), .Y(n12180) );
  INVX1_RVT U12311 ( .A(n12179), .Y(n12181) );
  INVX1_RVT U12312 ( .A(n11491), .Y(n12182) );
  INVX1_RVT U12313 ( .A(n12182), .Y(n12183) );
  INVX1_RVT U12314 ( .A(n1375), .Y(n12184) );
  INVX1_RVT U12315 ( .A(n12184), .Y(n12185) );
  INVX1_RVT U12316 ( .A(n12184), .Y(n12186) );
  INVX1_RVT U12317 ( .A(n1309), .Y(n12187) );
  INVX1_RVT U12318 ( .A(n12187), .Y(n12188) );
  INVX1_RVT U12319 ( .A(n12187), .Y(n12189) );
  INVX1_RVT U12320 ( .A(n6183), .Y(n12190) );
  INVX1_RVT U12321 ( .A(n12190), .Y(n12191) );
  INVX1_RVT U12322 ( .A(n12190), .Y(n12192) );
  INVX1_RVT U12323 ( .A(n1350), .Y(n12193) );
  INVX1_RVT U12324 ( .A(n12193), .Y(n12194) );
  XOR2X1_RVT U12325 ( .A1(key[100]), .A2(state[100]), .Y(n12195) );
  XOR2X1_RVT U12326 ( .A1(key[100]), .A2(state[100]), .Y(n12196) );
  INVX1_RVT U12327 ( .A(n1341), .Y(n12197) );
  INVX1_RVT U12328 ( .A(n12197), .Y(n12198) );
  INVX1_RVT U12329 ( .A(n12197), .Y(n12199) );
  INVX1_RVT U12330 ( .A(n1307), .Y(n12200) );
  INVX1_RVT U12331 ( .A(n12200), .Y(n12201) );
  INVX1_RVT U12332 ( .A(n1300), .Y(n12202) );
  INVX1_RVT U12333 ( .A(n12202), .Y(n12203) );
  INVX1_RVT U12334 ( .A(n12202), .Y(n12204) );
  INVX1_RVT U12335 ( .A(n1388), .Y(n12205) );
  INVX1_RVT U12336 ( .A(n12205), .Y(n12206) );
  INVX1_RVT U12337 ( .A(n6145), .Y(n12207) );
  INVX1_RVT U12338 ( .A(n12207), .Y(n12208) );
  INVX1_RVT U12339 ( .A(n12207), .Y(n12209) );
  INVX1_RVT U12340 ( .A(n1356), .Y(n12210) );
  INVX1_RVT U12341 ( .A(n12210), .Y(n12211) );
  INVX1_RVT U12342 ( .A(n12210), .Y(n12212) );
  INVX1_RVT U12343 ( .A(n10565), .Y(n12213) );
  INVX1_RVT U12344 ( .A(n12213), .Y(n12214) );
  XOR2X1_RVT U12345 ( .A1(key[81]), .A2(state[81]), .Y(n12215) );
  XOR2X1_RVT U12346 ( .A1(key[81]), .A2(state[81]), .Y(n12216) );
  INVX1_RVT U12347 ( .A(n10571), .Y(n12217) );
  INVX1_RVT U12348 ( .A(n12217), .Y(n12218) );
  INVX1_RVT U12349 ( .A(n12217), .Y(n12219) );
  INVX1_RVT U12350 ( .A(n10556), .Y(n12220) );
  INVX1_RVT U12351 ( .A(n12220), .Y(n12221) );
  INVX1_RVT U12352 ( .A(n10570), .Y(n12222) );
  INVX1_RVT U12353 ( .A(n12222), .Y(n12223) );
  INVX1_RVT U12354 ( .A(n10630), .Y(n12224) );
  INVX1_RVT U12355 ( .A(n12224), .Y(n12225) );
  INVX1_RVT U12356 ( .A(n12224), .Y(n12226) );
  INVX1_RVT U12357 ( .A(n12224), .Y(n12227) );
  INVX1_RVT U12358 ( .A(n10594), .Y(n12228) );
  INVX1_RVT U12359 ( .A(n12228), .Y(n12229) );
  INVX1_RVT U12360 ( .A(n12228), .Y(n12230) );
  INVX1_RVT U12361 ( .A(n12844), .Y(n12231) );
  INVX1_RVT U12362 ( .A(n12845), .Y(n12232) );
  INVX1_RVT U12363 ( .A(n10573), .Y(n12233) );
  INVX1_RVT U12364 ( .A(n12233), .Y(n12234) );
  INVX1_RVT U12365 ( .A(n10552), .Y(n12235) );
  INVX1_RVT U12366 ( .A(n12235), .Y(n12236) );
  INVX1_RVT U12367 ( .A(n12235), .Y(n12237) );
  INVX1_RVT U12368 ( .A(n10531), .Y(n12238) );
  INVX1_RVT U12369 ( .A(n12238), .Y(n12239) );
  INVX1_RVT U12370 ( .A(n12238), .Y(n12240) );
  INVX1_RVT U12371 ( .A(n10587), .Y(n12241) );
  INVX1_RVT U12372 ( .A(n12241), .Y(n12242) );
  INVX1_RVT U12373 ( .A(n12241), .Y(n12243) );
  INVX1_RVT U12374 ( .A(n10670), .Y(n12244) );
  INVX1_RVT U12375 ( .A(n12244), .Y(n12245) );
  INVX1_RVT U12376 ( .A(n9746), .Y(n12246) );
  INVX1_RVT U12377 ( .A(n12246), .Y(n12247) );
  XOR2X1_RVT U12378 ( .A1(key[89]), .A2(state[89]), .Y(n12248) );
  XOR2X1_RVT U12379 ( .A1(key[89]), .A2(state[89]), .Y(n12249) );
  INVX1_RVT U12380 ( .A(n9752), .Y(n12250) );
  INVX1_RVT U12381 ( .A(n12250), .Y(n12251) );
  INVX1_RVT U12382 ( .A(n12250), .Y(n12252) );
  INVX1_RVT U12383 ( .A(n9737), .Y(n12253) );
  INVX1_RVT U12384 ( .A(n12253), .Y(n12254) );
  INVX1_RVT U12385 ( .A(n9751), .Y(n12255) );
  INVX1_RVT U12386 ( .A(n12255), .Y(n12256) );
  INVX1_RVT U12387 ( .A(n9811), .Y(n12257) );
  INVX1_RVT U12388 ( .A(n12257), .Y(n12258) );
  INVX1_RVT U12389 ( .A(n12257), .Y(n12259) );
  INVX1_RVT U12390 ( .A(n12257), .Y(n12260) );
  INVX1_RVT U12391 ( .A(n9775), .Y(n12261) );
  INVX1_RVT U12392 ( .A(n12261), .Y(n12262) );
  INVX1_RVT U12393 ( .A(n12261), .Y(n12263) );
  INVX1_RVT U12394 ( .A(n12860), .Y(n12264) );
  INVX1_RVT U12395 ( .A(n12861), .Y(n12265) );
  INVX1_RVT U12396 ( .A(n9754), .Y(n12266) );
  INVX1_RVT U12397 ( .A(n12266), .Y(n12267) );
  INVX1_RVT U12398 ( .A(n9733), .Y(n12268) );
  INVX1_RVT U12399 ( .A(n12268), .Y(n12269) );
  INVX1_RVT U12400 ( .A(n12268), .Y(n12270) );
  INVX1_RVT U12401 ( .A(n9712), .Y(n12271) );
  INVX1_RVT U12402 ( .A(n12271), .Y(n12272) );
  INVX1_RVT U12403 ( .A(n12271), .Y(n12273) );
  INVX1_RVT U12404 ( .A(n9768), .Y(n12274) );
  INVX1_RVT U12405 ( .A(n12274), .Y(n12275) );
  INVX1_RVT U12406 ( .A(n12274), .Y(n12276) );
  INVX1_RVT U12407 ( .A(n9851), .Y(n12277) );
  INVX1_RVT U12408 ( .A(n12277), .Y(n12278) );
  INVX1_RVT U12409 ( .A(n9006), .Y(n12279) );
  INVX1_RVT U12410 ( .A(n12279), .Y(n12280) );
  XOR2X1_RVT U12411 ( .A1(key[33]), .A2(state[33]), .Y(n12281) );
  XOR2X1_RVT U12412 ( .A1(key[33]), .A2(state[33]), .Y(n12282) );
  INVX1_RVT U12413 ( .A(n9012), .Y(n12283) );
  INVX1_RVT U12414 ( .A(n12283), .Y(n12284) );
  INVX1_RVT U12415 ( .A(n12283), .Y(n12285) );
  INVX1_RVT U12416 ( .A(n8997), .Y(n12286) );
  INVX1_RVT U12417 ( .A(n12286), .Y(n12287) );
  INVX1_RVT U12418 ( .A(n9011), .Y(n12288) );
  INVX1_RVT U12419 ( .A(n12288), .Y(n12289) );
  INVX1_RVT U12420 ( .A(n9071), .Y(n12290) );
  INVX1_RVT U12421 ( .A(n12290), .Y(n12291) );
  INVX1_RVT U12422 ( .A(n12290), .Y(n12292) );
  INVX1_RVT U12423 ( .A(n12290), .Y(n12293) );
  INVX1_RVT U12424 ( .A(n9035), .Y(n12294) );
  INVX1_RVT U12425 ( .A(n12294), .Y(n12295) );
  INVX1_RVT U12426 ( .A(n12294), .Y(n12296) );
  INVX1_RVT U12427 ( .A(n12748), .Y(n12297) );
  INVX1_RVT U12428 ( .A(n12749), .Y(n12298) );
  INVX1_RVT U12429 ( .A(n9014), .Y(n12299) );
  INVX1_RVT U12430 ( .A(n12299), .Y(n12300) );
  INVX1_RVT U12431 ( .A(n8993), .Y(n12301) );
  INVX1_RVT U12432 ( .A(n12301), .Y(n12302) );
  INVX1_RVT U12433 ( .A(n12301), .Y(n12303) );
  INVX1_RVT U12434 ( .A(n8972), .Y(n12304) );
  INVX1_RVT U12435 ( .A(n12304), .Y(n12305) );
  INVX1_RVT U12436 ( .A(n12304), .Y(n12306) );
  INVX1_RVT U12437 ( .A(n9028), .Y(n12307) );
  INVX1_RVT U12438 ( .A(n12307), .Y(n12308) );
  INVX1_RVT U12439 ( .A(n12307), .Y(n12309) );
  INVX1_RVT U12440 ( .A(n9111), .Y(n12310) );
  INVX1_RVT U12441 ( .A(n12310), .Y(n12311) );
  INVX1_RVT U12442 ( .A(n8182), .Y(n12312) );
  INVX1_RVT U12443 ( .A(n12312), .Y(n12313) );
  XOR2X1_RVT U12444 ( .A1(key[41]), .A2(state[41]), .Y(n12314) );
  XOR2X1_RVT U12445 ( .A1(key[41]), .A2(state[41]), .Y(n12315) );
  INVX1_RVT U12446 ( .A(n8188), .Y(n12316) );
  INVX1_RVT U12447 ( .A(n12316), .Y(n12317) );
  INVX1_RVT U12448 ( .A(n12316), .Y(n12318) );
  INVX1_RVT U12449 ( .A(n8173), .Y(n12319) );
  INVX1_RVT U12450 ( .A(n12319), .Y(n12320) );
  INVX1_RVT U12451 ( .A(n8187), .Y(n12321) );
  INVX1_RVT U12452 ( .A(n12321), .Y(n12322) );
  INVX1_RVT U12453 ( .A(n8247), .Y(n12323) );
  INVX1_RVT U12454 ( .A(n12323), .Y(n12324) );
  INVX1_RVT U12455 ( .A(n12323), .Y(n12325) );
  INVX1_RVT U12456 ( .A(n12323), .Y(n12326) );
  INVX1_RVT U12457 ( .A(n8211), .Y(n12327) );
  INVX1_RVT U12458 ( .A(n12327), .Y(n12328) );
  INVX1_RVT U12459 ( .A(n12327), .Y(n12329) );
  INVX1_RVT U12460 ( .A(n12764), .Y(n12330) );
  INVX1_RVT U12461 ( .A(n12765), .Y(n12331) );
  INVX1_RVT U12462 ( .A(n8190), .Y(n12332) );
  INVX1_RVT U12463 ( .A(n12332), .Y(n12333) );
  INVX1_RVT U12464 ( .A(n8169), .Y(n12334) );
  INVX1_RVT U12465 ( .A(n12334), .Y(n12335) );
  INVX1_RVT U12466 ( .A(n12334), .Y(n12336) );
  INVX1_RVT U12467 ( .A(n8148), .Y(n12337) );
  INVX1_RVT U12468 ( .A(n12337), .Y(n12338) );
  INVX1_RVT U12469 ( .A(n12337), .Y(n12339) );
  INVX1_RVT U12470 ( .A(n8204), .Y(n12340) );
  INVX1_RVT U12471 ( .A(n12340), .Y(n12341) );
  INVX1_RVT U12472 ( .A(n12340), .Y(n12342) );
  INVX1_RVT U12473 ( .A(n8287), .Y(n12343) );
  INVX1_RVT U12474 ( .A(n12343), .Y(n12344) );
  INVX1_RVT U12475 ( .A(n7351), .Y(n12345) );
  INVX1_RVT U12476 ( .A(n12345), .Y(n12346) );
  XOR2X1_RVT U12477 ( .A1(key[49]), .A2(state[49]), .Y(n12347) );
  XOR2X1_RVT U12478 ( .A1(key[49]), .A2(state[49]), .Y(n12348) );
  INVX1_RVT U12479 ( .A(n7357), .Y(n12349) );
  INVX1_RVT U12480 ( .A(n12349), .Y(n12350) );
  INVX1_RVT U12481 ( .A(n12349), .Y(n12351) );
  INVX1_RVT U12482 ( .A(n7342), .Y(n12352) );
  INVX1_RVT U12483 ( .A(n12352), .Y(n12353) );
  INVX1_RVT U12484 ( .A(n7356), .Y(n12354) );
  INVX1_RVT U12485 ( .A(n12354), .Y(n12355) );
  INVX1_RVT U12486 ( .A(n7416), .Y(n12356) );
  INVX1_RVT U12487 ( .A(n12356), .Y(n12357) );
  INVX1_RVT U12488 ( .A(n12356), .Y(n12358) );
  INVX1_RVT U12489 ( .A(n12356), .Y(n12359) );
  INVX1_RVT U12490 ( .A(n7380), .Y(n12360) );
  INVX1_RVT U12491 ( .A(n12360), .Y(n12361) );
  INVX1_RVT U12492 ( .A(n12360), .Y(n12362) );
  INVX1_RVT U12493 ( .A(n12780), .Y(n12363) );
  INVX1_RVT U12494 ( .A(n12781), .Y(n12364) );
  INVX1_RVT U12495 ( .A(n7359), .Y(n12365) );
  INVX1_RVT U12496 ( .A(n12365), .Y(n12366) );
  INVX1_RVT U12497 ( .A(n7338), .Y(n12367) );
  INVX1_RVT U12498 ( .A(n12367), .Y(n12368) );
  INVX1_RVT U12499 ( .A(n12367), .Y(n12369) );
  INVX1_RVT U12500 ( .A(n7317), .Y(n12370) );
  INVX1_RVT U12501 ( .A(n12370), .Y(n12371) );
  INVX1_RVT U12502 ( .A(n12370), .Y(n12372) );
  INVX1_RVT U12503 ( .A(n7373), .Y(n12373) );
  INVX1_RVT U12504 ( .A(n12373), .Y(n12374) );
  INVX1_RVT U12505 ( .A(n12373), .Y(n12375) );
  INVX1_RVT U12506 ( .A(n7456), .Y(n12376) );
  INVX1_RVT U12507 ( .A(n12376), .Y(n12377) );
  INVX1_RVT U12508 ( .A(n6512), .Y(n12378) );
  INVX1_RVT U12509 ( .A(n12378), .Y(n12379) );
  XOR2X1_RVT U12510 ( .A1(key[57]), .A2(state[57]), .Y(n12380) );
  XOR2X1_RVT U12511 ( .A1(key[57]), .A2(state[57]), .Y(n12381) );
  INVX1_RVT U12512 ( .A(n6518), .Y(n12382) );
  INVX1_RVT U12513 ( .A(n12382), .Y(n12383) );
  INVX1_RVT U12514 ( .A(n12382), .Y(n12384) );
  INVX1_RVT U12515 ( .A(n6503), .Y(n12385) );
  INVX1_RVT U12516 ( .A(n12385), .Y(n12386) );
  INVX1_RVT U12517 ( .A(n6517), .Y(n12387) );
  INVX1_RVT U12518 ( .A(n12387), .Y(n12388) );
  INVX1_RVT U12519 ( .A(n6577), .Y(n12389) );
  INVX1_RVT U12520 ( .A(n12389), .Y(n12390) );
  INVX1_RVT U12521 ( .A(n12389), .Y(n12391) );
  INVX1_RVT U12522 ( .A(n12389), .Y(n12392) );
  INVX1_RVT U12523 ( .A(n6541), .Y(n12393) );
  INVX1_RVT U12524 ( .A(n12393), .Y(n12394) );
  INVX1_RVT U12525 ( .A(n12393), .Y(n12395) );
  INVX1_RVT U12526 ( .A(n12796), .Y(n12396) );
  INVX1_RVT U12527 ( .A(n12797), .Y(n12397) );
  INVX1_RVT U12528 ( .A(n6520), .Y(n12398) );
  INVX1_RVT U12529 ( .A(n12398), .Y(n12399) );
  INVX1_RVT U12530 ( .A(n6499), .Y(n12400) );
  INVX1_RVT U12531 ( .A(n12400), .Y(n12401) );
  INVX1_RVT U12532 ( .A(n12400), .Y(n12402) );
  INVX1_RVT U12533 ( .A(n6478), .Y(n12403) );
  INVX1_RVT U12534 ( .A(n12403), .Y(n12404) );
  INVX1_RVT U12535 ( .A(n12403), .Y(n12405) );
  INVX1_RVT U12536 ( .A(n6534), .Y(n12406) );
  INVX1_RVT U12537 ( .A(n12406), .Y(n12407) );
  INVX1_RVT U12538 ( .A(n12406), .Y(n12408) );
  INVX1_RVT U12539 ( .A(n6617), .Y(n12409) );
  INVX1_RVT U12540 ( .A(n12409), .Y(n12410) );
  INVX1_RVT U12541 ( .A(n5672), .Y(n12411) );
  INVX1_RVT U12542 ( .A(n12411), .Y(n12412) );
  XOR2X1_RVT U12543 ( .A1(key[1]), .A2(state[1]), .Y(n12413) );
  XOR2X1_RVT U12544 ( .A1(key[1]), .A2(state[1]), .Y(n12414) );
  INVX1_RVT U12545 ( .A(n5678), .Y(n12415) );
  INVX1_RVT U12546 ( .A(n12415), .Y(n12416) );
  INVX1_RVT U12547 ( .A(n12415), .Y(n12417) );
  INVX1_RVT U12548 ( .A(n5663), .Y(n12418) );
  INVX1_RVT U12549 ( .A(n12418), .Y(n12419) );
  INVX1_RVT U12550 ( .A(n5677), .Y(n12420) );
  INVX1_RVT U12551 ( .A(n12420), .Y(n12421) );
  INVX1_RVT U12552 ( .A(n5737), .Y(n12422) );
  INVX1_RVT U12553 ( .A(n12422), .Y(n12423) );
  INVX1_RVT U12554 ( .A(n12422), .Y(n12424) );
  INVX1_RVT U12555 ( .A(n12422), .Y(n12425) );
  INVX1_RVT U12556 ( .A(n5701), .Y(n12426) );
  INVX1_RVT U12557 ( .A(n12426), .Y(n12427) );
  INVX1_RVT U12558 ( .A(n12426), .Y(n12428) );
  INVX1_RVT U12559 ( .A(n12684), .Y(n12429) );
  INVX1_RVT U12560 ( .A(n12685), .Y(n12430) );
  INVX1_RVT U12561 ( .A(n5680), .Y(n12431) );
  INVX1_RVT U12562 ( .A(n12431), .Y(n12432) );
  INVX1_RVT U12563 ( .A(n5659), .Y(n12433) );
  INVX1_RVT U12564 ( .A(n12433), .Y(n12434) );
  INVX1_RVT U12565 ( .A(n12433), .Y(n12435) );
  INVX1_RVT U12566 ( .A(n5638), .Y(n12436) );
  INVX1_RVT U12567 ( .A(n12436), .Y(n12437) );
  INVX1_RVT U12568 ( .A(n12436), .Y(n12438) );
  INVX1_RVT U12569 ( .A(n5694), .Y(n12439) );
  INVX1_RVT U12570 ( .A(n12439), .Y(n12440) );
  INVX1_RVT U12571 ( .A(n12439), .Y(n12441) );
  INVX1_RVT U12572 ( .A(n5777), .Y(n12442) );
  INVX1_RVT U12573 ( .A(n12442), .Y(n12443) );
  INVX1_RVT U12574 ( .A(n4849), .Y(n12444) );
  INVX1_RVT U12575 ( .A(n12444), .Y(n12445) );
  XOR2X1_RVT U12576 ( .A1(key[9]), .A2(state[9]), .Y(n12446) );
  XOR2X1_RVT U12577 ( .A1(key[9]), .A2(state[9]), .Y(n12447) );
  INVX1_RVT U12578 ( .A(n4855), .Y(n12448) );
  INVX1_RVT U12579 ( .A(n12448), .Y(n12449) );
  INVX1_RVT U12580 ( .A(n12448), .Y(n12450) );
  INVX1_RVT U12581 ( .A(n4840), .Y(n12451) );
  INVX1_RVT U12582 ( .A(n12451), .Y(n12452) );
  INVX1_RVT U12583 ( .A(n4854), .Y(n12453) );
  INVX1_RVT U12584 ( .A(n12453), .Y(n12454) );
  INVX1_RVT U12585 ( .A(n4914), .Y(n12455) );
  INVX1_RVT U12586 ( .A(n12455), .Y(n12456) );
  INVX1_RVT U12587 ( .A(n12455), .Y(n12457) );
  INVX1_RVT U12588 ( .A(n12455), .Y(n12458) );
  INVX1_RVT U12589 ( .A(n4878), .Y(n12459) );
  INVX1_RVT U12590 ( .A(n12459), .Y(n12460) );
  INVX1_RVT U12591 ( .A(n12459), .Y(n12461) );
  INVX1_RVT U12592 ( .A(n12700), .Y(n12462) );
  INVX1_RVT U12593 ( .A(n12701), .Y(n12463) );
  INVX1_RVT U12594 ( .A(n4857), .Y(n12464) );
  INVX1_RVT U12595 ( .A(n12464), .Y(n12465) );
  INVX1_RVT U12596 ( .A(n4836), .Y(n12466) );
  INVX1_RVT U12597 ( .A(n12466), .Y(n12467) );
  INVX1_RVT U12598 ( .A(n12466), .Y(n12468) );
  INVX1_RVT U12599 ( .A(n4815), .Y(n12469) );
  INVX1_RVT U12600 ( .A(n12469), .Y(n12470) );
  INVX1_RVT U12601 ( .A(n12469), .Y(n12471) );
  INVX1_RVT U12602 ( .A(n4871), .Y(n12472) );
  INVX1_RVT U12603 ( .A(n12472), .Y(n12473) );
  INVX1_RVT U12604 ( .A(n12472), .Y(n12474) );
  INVX1_RVT U12605 ( .A(n4954), .Y(n12475) );
  INVX1_RVT U12606 ( .A(n12475), .Y(n12476) );
  INVX1_RVT U12607 ( .A(n2712), .Y(n12477) );
  INVX1_RVT U12608 ( .A(n12477), .Y(n12478) );
  XOR2X1_RVT U12609 ( .A1(key[105]), .A2(state[105]), .Y(n12479) );
  XOR2X1_RVT U12610 ( .A1(key[105]), .A2(state[105]), .Y(n12480) );
  INVX1_RVT U12611 ( .A(n2718), .Y(n12481) );
  INVX1_RVT U12612 ( .A(n12481), .Y(n12482) );
  INVX1_RVT U12613 ( .A(n12481), .Y(n12483) );
  INVX1_RVT U12614 ( .A(n2703), .Y(n12484) );
  INVX1_RVT U12615 ( .A(n12484), .Y(n12485) );
  INVX1_RVT U12616 ( .A(n2717), .Y(n12486) );
  INVX1_RVT U12617 ( .A(n12486), .Y(n12487) );
  INVX1_RVT U12618 ( .A(n2777), .Y(n12488) );
  INVX1_RVT U12619 ( .A(n12488), .Y(n12489) );
  INVX1_RVT U12620 ( .A(n12488), .Y(n12490) );
  INVX1_RVT U12621 ( .A(n12488), .Y(n12491) );
  INVX1_RVT U12622 ( .A(n2741), .Y(n12492) );
  INVX1_RVT U12623 ( .A(n12492), .Y(n12493) );
  INVX1_RVT U12624 ( .A(n12492), .Y(n12494) );
  INVX1_RVT U12625 ( .A(n12887), .Y(n12495) );
  INVX1_RVT U12626 ( .A(n12888), .Y(n12496) );
  INVX1_RVT U12627 ( .A(n2720), .Y(n12497) );
  INVX1_RVT U12628 ( .A(n12497), .Y(n12498) );
  INVX1_RVT U12629 ( .A(n2699), .Y(n12499) );
  INVX1_RVT U12630 ( .A(n12499), .Y(n12500) );
  INVX1_RVT U12631 ( .A(n12499), .Y(n12501) );
  INVX1_RVT U12632 ( .A(n2678), .Y(n12502) );
  INVX1_RVT U12633 ( .A(n12502), .Y(n12503) );
  INVX1_RVT U12634 ( .A(n12502), .Y(n12504) );
  INVX1_RVT U12635 ( .A(n2734), .Y(n12505) );
  INVX1_RVT U12636 ( .A(n12505), .Y(n12506) );
  INVX1_RVT U12637 ( .A(n12505), .Y(n12507) );
  INVX1_RVT U12638 ( .A(n2817), .Y(n12508) );
  INVX1_RVT U12639 ( .A(n12508), .Y(n12509) );
  INVX1_RVT U12640 ( .A(n4109), .Y(n12510) );
  INVX1_RVT U12641 ( .A(n12510), .Y(n12511) );
  XOR2X1_RVT U12642 ( .A1(key[17]), .A2(state[17]), .Y(n12512) );
  XOR2X1_RVT U12643 ( .A1(key[17]), .A2(state[17]), .Y(n12513) );
  INVX1_RVT U12644 ( .A(n4115), .Y(n12514) );
  INVX1_RVT U12645 ( .A(n12514), .Y(n12515) );
  INVX1_RVT U12646 ( .A(n12514), .Y(n12516) );
  INVX1_RVT U12647 ( .A(n4100), .Y(n12517) );
  INVX1_RVT U12648 ( .A(n12517), .Y(n12518) );
  INVX1_RVT U12649 ( .A(n4114), .Y(n12519) );
  INVX1_RVT U12650 ( .A(n12519), .Y(n12520) );
  INVX1_RVT U12651 ( .A(n4174), .Y(n12521) );
  INVX1_RVT U12652 ( .A(n12521), .Y(n12522) );
  INVX1_RVT U12653 ( .A(n12521), .Y(n12523) );
  INVX1_RVT U12654 ( .A(n12521), .Y(n12524) );
  INVX1_RVT U12655 ( .A(n4138), .Y(n12525) );
  INVX1_RVT U12656 ( .A(n12525), .Y(n12526) );
  INVX1_RVT U12657 ( .A(n12525), .Y(n12527) );
  INVX1_RVT U12658 ( .A(n12716), .Y(n12528) );
  INVX1_RVT U12659 ( .A(n12717), .Y(n12529) );
  INVX1_RVT U12660 ( .A(n4117), .Y(n12530) );
  INVX1_RVT U12661 ( .A(n12530), .Y(n12531) );
  INVX1_RVT U12662 ( .A(n4096), .Y(n12532) );
  INVX1_RVT U12663 ( .A(n12532), .Y(n12533) );
  INVX1_RVT U12664 ( .A(n12532), .Y(n12534) );
  INVX1_RVT U12665 ( .A(n4075), .Y(n12535) );
  INVX1_RVT U12666 ( .A(n12535), .Y(n12536) );
  INVX1_RVT U12667 ( .A(n12535), .Y(n12537) );
  INVX1_RVT U12668 ( .A(n4131), .Y(n12538) );
  INVX1_RVT U12669 ( .A(n12538), .Y(n12539) );
  INVX1_RVT U12670 ( .A(n12538), .Y(n12540) );
  INVX1_RVT U12671 ( .A(n4214), .Y(n12541) );
  INVX1_RVT U12672 ( .A(n12541), .Y(n12542) );
  INVX1_RVT U12673 ( .A(n3292), .Y(n12543) );
  INVX1_RVT U12674 ( .A(n12543), .Y(n12544) );
  XOR2X1_RVT U12675 ( .A1(key[25]), .A2(state[25]), .Y(n12545) );
  XOR2X1_RVT U12676 ( .A1(key[25]), .A2(state[25]), .Y(n12546) );
  INVX1_RVT U12677 ( .A(n3298), .Y(n12547) );
  INVX1_RVT U12678 ( .A(n12547), .Y(n12548) );
  INVX1_RVT U12679 ( .A(n12547), .Y(n12549) );
  INVX1_RVT U12680 ( .A(n3283), .Y(n12550) );
  INVX1_RVT U12681 ( .A(n12550), .Y(n12551) );
  INVX1_RVT U12682 ( .A(n3297), .Y(n12552) );
  INVX1_RVT U12683 ( .A(n12552), .Y(n12553) );
  INVX1_RVT U12684 ( .A(n3357), .Y(n12554) );
  INVX1_RVT U12685 ( .A(n12554), .Y(n12555) );
  INVX1_RVT U12686 ( .A(n12554), .Y(n12556) );
  INVX1_RVT U12687 ( .A(n12554), .Y(n12557) );
  INVX1_RVT U12688 ( .A(n3321), .Y(n12558) );
  INVX1_RVT U12689 ( .A(n12558), .Y(n12559) );
  INVX1_RVT U12690 ( .A(n12558), .Y(n12560) );
  INVX1_RVT U12691 ( .A(n12732), .Y(n12561) );
  INVX1_RVT U12692 ( .A(n12733), .Y(n12562) );
  INVX1_RVT U12693 ( .A(n3300), .Y(n12563) );
  INVX1_RVT U12694 ( .A(n12563), .Y(n12564) );
  INVX1_RVT U12695 ( .A(n3279), .Y(n12565) );
  INVX1_RVT U12696 ( .A(n12565), .Y(n12566) );
  INVX1_RVT U12697 ( .A(n12565), .Y(n12567) );
  INVX1_RVT U12698 ( .A(n3258), .Y(n12568) );
  INVX1_RVT U12699 ( .A(n12568), .Y(n12569) );
  INVX1_RVT U12700 ( .A(n12568), .Y(n12570) );
  INVX1_RVT U12701 ( .A(n3314), .Y(n12571) );
  INVX1_RVT U12702 ( .A(n12571), .Y(n12572) );
  INVX1_RVT U12703 ( .A(n12571), .Y(n12573) );
  INVX1_RVT U12704 ( .A(n3397), .Y(n12574) );
  INVX1_RVT U12705 ( .A(n12574), .Y(n12575) );
  INVX1_RVT U12706 ( .A(n1972), .Y(n12576) );
  INVX1_RVT U12707 ( .A(n12576), .Y(n12577) );
  XOR2X1_RVT U12708 ( .A1(key[113]), .A2(state[113]), .Y(n12578) );
  XOR2X1_RVT U12709 ( .A1(key[113]), .A2(state[113]), .Y(n12579) );
  INVX1_RVT U12710 ( .A(n1978), .Y(n12580) );
  INVX1_RVT U12711 ( .A(n12580), .Y(n12581) );
  INVX1_RVT U12712 ( .A(n12580), .Y(n12582) );
  INVX1_RVT U12713 ( .A(n1963), .Y(n12583) );
  INVX1_RVT U12714 ( .A(n12583), .Y(n12584) );
  INVX1_RVT U12715 ( .A(n1977), .Y(n12585) );
  INVX1_RVT U12716 ( .A(n12585), .Y(n12586) );
  INVX1_RVT U12717 ( .A(n2037), .Y(n12587) );
  INVX1_RVT U12718 ( .A(n12587), .Y(n12588) );
  INVX1_RVT U12719 ( .A(n12587), .Y(n12589) );
  INVX1_RVT U12720 ( .A(n12587), .Y(n12590) );
  INVX1_RVT U12721 ( .A(n2001), .Y(n12591) );
  INVX1_RVT U12722 ( .A(n12591), .Y(n12592) );
  INVX1_RVT U12723 ( .A(n12591), .Y(n12593) );
  INVX1_RVT U12724 ( .A(n12903), .Y(n12594) );
  INVX1_RVT U12725 ( .A(n12904), .Y(n12595) );
  INVX1_RVT U12726 ( .A(n1980), .Y(n12596) );
  INVX1_RVT U12727 ( .A(n12596), .Y(n12597) );
  INVX1_RVT U12728 ( .A(n1959), .Y(n12598) );
  INVX1_RVT U12729 ( .A(n12598), .Y(n12599) );
  INVX1_RVT U12730 ( .A(n12598), .Y(n12600) );
  INVX1_RVT U12731 ( .A(n1938), .Y(n12601) );
  INVX1_RVT U12732 ( .A(n12601), .Y(n12602) );
  INVX1_RVT U12733 ( .A(n12601), .Y(n12603) );
  INVX1_RVT U12734 ( .A(n1994), .Y(n12604) );
  INVX1_RVT U12735 ( .A(n12604), .Y(n12605) );
  INVX1_RVT U12736 ( .A(n12604), .Y(n12606) );
  INVX1_RVT U12737 ( .A(n2077), .Y(n12607) );
  INVX1_RVT U12738 ( .A(n12607), .Y(n12608) );
  INVX1_RVT U12739 ( .A(n1113), .Y(n12609) );
  INVX1_RVT U12740 ( .A(n12609), .Y(n12610) );
  XOR2X1_RVT U12741 ( .A1(key[121]), .A2(state[121]), .Y(n12611) );
  XOR2X1_RVT U12742 ( .A1(key[121]), .A2(state[121]), .Y(n12612) );
  INVX1_RVT U12743 ( .A(n1119), .Y(n12613) );
  INVX1_RVT U12744 ( .A(n12613), .Y(n12614) );
  INVX1_RVT U12745 ( .A(n12613), .Y(n12615) );
  INVX1_RVT U12746 ( .A(n1104), .Y(n12616) );
  INVX1_RVT U12747 ( .A(n12616), .Y(n12617) );
  INVX1_RVT U12748 ( .A(n1118), .Y(n12618) );
  INVX1_RVT U12749 ( .A(n12618), .Y(n12619) );
  INVX1_RVT U12750 ( .A(n1178), .Y(n12620) );
  INVX1_RVT U12751 ( .A(n12620), .Y(n12621) );
  INVX1_RVT U12752 ( .A(n12620), .Y(n12622) );
  INVX1_RVT U12753 ( .A(n12620), .Y(n12623) );
  INVX1_RVT U12754 ( .A(n1142), .Y(n12624) );
  INVX1_RVT U12755 ( .A(n12624), .Y(n12625) );
  INVX1_RVT U12756 ( .A(n12624), .Y(n12626) );
  INVX1_RVT U12757 ( .A(n12919), .Y(n12627) );
  INVX1_RVT U12758 ( .A(n12920), .Y(n12628) );
  INVX1_RVT U12759 ( .A(n1121), .Y(n12629) );
  INVX1_RVT U12760 ( .A(n12629), .Y(n12630) );
  INVX1_RVT U12761 ( .A(n1100), .Y(n12631) );
  INVX1_RVT U12762 ( .A(n12631), .Y(n12632) );
  INVX1_RVT U12763 ( .A(n12631), .Y(n12633) );
  INVX1_RVT U12764 ( .A(n1079), .Y(n12634) );
  INVX1_RVT U12765 ( .A(n12634), .Y(n12635) );
  INVX1_RVT U12766 ( .A(n12634), .Y(n12636) );
  INVX1_RVT U12767 ( .A(n1135), .Y(n12637) );
  INVX1_RVT U12768 ( .A(n12637), .Y(n12638) );
  INVX1_RVT U12769 ( .A(n12637), .Y(n12639) );
  INVX1_RVT U12770 ( .A(n1218), .Y(n12640) );
  INVX1_RVT U12771 ( .A(n12640), .Y(n12641) );
  INVX1_RVT U12772 ( .A(n373), .Y(n12642) );
  INVX1_RVT U12773 ( .A(n12642), .Y(n12643) );
  XOR2X1_RVT U12774 ( .A1(key[65]), .A2(state[65]), .Y(n12644) );
  XOR2X1_RVT U12775 ( .A1(key[65]), .A2(state[65]), .Y(n12645) );
  INVX1_RVT U12776 ( .A(n379), .Y(n12646) );
  INVX1_RVT U12777 ( .A(n12646), .Y(n12647) );
  INVX1_RVT U12778 ( .A(n12646), .Y(n12648) );
  INVX1_RVT U12779 ( .A(n364), .Y(n12649) );
  INVX1_RVT U12780 ( .A(n12649), .Y(n12650) );
  INVX1_RVT U12781 ( .A(n378), .Y(n12651) );
  INVX1_RVT U12782 ( .A(n12651), .Y(n12652) );
  INVX1_RVT U12783 ( .A(n438), .Y(n12653) );
  INVX1_RVT U12784 ( .A(n12653), .Y(n12654) );
  INVX1_RVT U12785 ( .A(n12653), .Y(n12655) );
  INVX1_RVT U12786 ( .A(n12653), .Y(n12656) );
  INVX1_RVT U12787 ( .A(n402), .Y(n12657) );
  INVX1_RVT U12788 ( .A(n12657), .Y(n12658) );
  INVX1_RVT U12789 ( .A(n12657), .Y(n12659) );
  INVX1_RVT U12790 ( .A(n12812), .Y(n12660) );
  INVX1_RVT U12791 ( .A(n12813), .Y(n12661) );
  INVX1_RVT U12792 ( .A(n381), .Y(n12662) );
  INVX1_RVT U12793 ( .A(n12662), .Y(n12663) );
  INVX1_RVT U12794 ( .A(n360), .Y(n12664) );
  INVX1_RVT U12795 ( .A(n12664), .Y(n12665) );
  INVX1_RVT U12796 ( .A(n12664), .Y(n12666) );
  INVX1_RVT U12797 ( .A(n339), .Y(n12667) );
  INVX1_RVT U12798 ( .A(n12667), .Y(n12668) );
  INVX1_RVT U12799 ( .A(n12667), .Y(n12669) );
  INVX1_RVT U12800 ( .A(n395), .Y(n12670) );
  INVX1_RVT U12801 ( .A(n12670), .Y(n12671) );
  INVX1_RVT U12802 ( .A(n12670), .Y(n12672) );
  INVX1_RVT U12803 ( .A(n478), .Y(n12673) );
  INVX1_RVT U12804 ( .A(n12673), .Y(n12674) );
  INVX1_RVT U12805 ( .A(n12416), .Y(n12675) );
  INVX1_RVT U12806 ( .A(n5678), .Y(n12676) );
  INVX1_RVT U12807 ( .A(n12414), .Y(n12677) );
  INVX1_RVT U12808 ( .A(n12414), .Y(n12678) );
  INVX1_RVT U12809 ( .A(n5803), .Y(n12679) );
  INVX1_RVT U12810 ( .A(n5803), .Y(n12680) );
  INVX1_RVT U12811 ( .A(n12425), .Y(n12681) );
  INVX1_RVT U12812 ( .A(n12423), .Y(n12682) );
  INVX1_RVT U12813 ( .A(n12424), .Y(n12683) );
  INVX1_RVT U12814 ( .A(n5655), .Y(n12684) );
  INVX1_RVT U12815 ( .A(n5655), .Y(n12685) );
  INVX1_RVT U12816 ( .A(n5752), .Y(n12686) );
  INVX1_RVT U12817 ( .A(n5752), .Y(n12687) );
  INVX1_RVT U12818 ( .A(n5699), .Y(n12688) );
  INVX1_RVT U12819 ( .A(n5699), .Y(n12689) );
  INVX1_RVT U12820 ( .A(n12412), .Y(n12690) );
  INVX1_RVT U12821 ( .A(n12449), .Y(n12691) );
  INVX1_RVT U12822 ( .A(n4855), .Y(n12692) );
  INVX1_RVT U12823 ( .A(n12447), .Y(n12693) );
  INVX1_RVT U12824 ( .A(n12447), .Y(n12694) );
  INVX1_RVT U12825 ( .A(n4980), .Y(n12695) );
  INVX1_RVT U12826 ( .A(n4980), .Y(n12696) );
  INVX1_RVT U12827 ( .A(n12458), .Y(n12697) );
  INVX1_RVT U12828 ( .A(n12456), .Y(n12698) );
  INVX1_RVT U12829 ( .A(n12457), .Y(n12699) );
  INVX1_RVT U12830 ( .A(n4832), .Y(n12700) );
  INVX1_RVT U12831 ( .A(n4832), .Y(n12701) );
  INVX1_RVT U12832 ( .A(n4929), .Y(n12702) );
  INVX1_RVT U12833 ( .A(n4929), .Y(n12703) );
  INVX1_RVT U12834 ( .A(n4876), .Y(n12704) );
  INVX1_RVT U12835 ( .A(n4876), .Y(n12705) );
  INVX1_RVT U12836 ( .A(n12445), .Y(n12706) );
  INVX1_RVT U12837 ( .A(n12515), .Y(n12707) );
  INVX1_RVT U12838 ( .A(n4115), .Y(n12708) );
  INVX1_RVT U12839 ( .A(n12513), .Y(n12709) );
  INVX1_RVT U12840 ( .A(n12513), .Y(n12710) );
  INVX1_RVT U12841 ( .A(n4240), .Y(n12711) );
  INVX1_RVT U12842 ( .A(n4240), .Y(n12712) );
  INVX1_RVT U12843 ( .A(n12524), .Y(n12713) );
  INVX1_RVT U12844 ( .A(n12522), .Y(n12714) );
  INVX1_RVT U12845 ( .A(n12523), .Y(n12715) );
  INVX1_RVT U12846 ( .A(n4092), .Y(n12716) );
  INVX1_RVT U12847 ( .A(n4092), .Y(n12717) );
  INVX1_RVT U12848 ( .A(n4189), .Y(n12718) );
  INVX1_RVT U12849 ( .A(n4189), .Y(n12719) );
  INVX1_RVT U12850 ( .A(n4136), .Y(n12720) );
  INVX1_RVT U12851 ( .A(n4136), .Y(n12721) );
  INVX1_RVT U12852 ( .A(n12511), .Y(n12722) );
  INVX1_RVT U12853 ( .A(n12548), .Y(n12723) );
  INVX1_RVT U12854 ( .A(n3298), .Y(n12724) );
  INVX1_RVT U12855 ( .A(n12546), .Y(n12725) );
  INVX1_RVT U12856 ( .A(n12546), .Y(n12726) );
  INVX1_RVT U12857 ( .A(n3423), .Y(n12727) );
  INVX1_RVT U12858 ( .A(n3423), .Y(n12728) );
  INVX1_RVT U12859 ( .A(n12557), .Y(n12729) );
  INVX1_RVT U12860 ( .A(n12555), .Y(n12730) );
  INVX1_RVT U12861 ( .A(n12556), .Y(n12731) );
  INVX1_RVT U12862 ( .A(n3275), .Y(n12732) );
  INVX1_RVT U12863 ( .A(n3275), .Y(n12733) );
  INVX1_RVT U12864 ( .A(n3372), .Y(n12734) );
  INVX1_RVT U12865 ( .A(n3372), .Y(n12735) );
  INVX1_RVT U12866 ( .A(n3319), .Y(n12736) );
  INVX1_RVT U12867 ( .A(n3319), .Y(n12737) );
  INVX1_RVT U12868 ( .A(n12544), .Y(n12738) );
  INVX1_RVT U12869 ( .A(n12284), .Y(n12739) );
  INVX1_RVT U12870 ( .A(n9012), .Y(n12740) );
  INVX1_RVT U12871 ( .A(n12282), .Y(n12741) );
  INVX1_RVT U12872 ( .A(n12282), .Y(n12742) );
  INVX1_RVT U12873 ( .A(n9137), .Y(n12743) );
  INVX1_RVT U12874 ( .A(n9137), .Y(n12744) );
  INVX1_RVT U12875 ( .A(n12293), .Y(n12745) );
  INVX1_RVT U12876 ( .A(n12291), .Y(n12746) );
  INVX1_RVT U12877 ( .A(n12292), .Y(n12747) );
  INVX1_RVT U12878 ( .A(n8989), .Y(n12748) );
  INVX1_RVT U12879 ( .A(n8989), .Y(n12749) );
  INVX1_RVT U12880 ( .A(n9086), .Y(n12750) );
  INVX1_RVT U12881 ( .A(n9086), .Y(n12751) );
  INVX1_RVT U12882 ( .A(n9033), .Y(n12752) );
  INVX1_RVT U12883 ( .A(n9033), .Y(n12753) );
  INVX1_RVT U12884 ( .A(n12280), .Y(n12754) );
  INVX1_RVT U12885 ( .A(n12317), .Y(n12755) );
  INVX1_RVT U12886 ( .A(n8188), .Y(n12756) );
  INVX1_RVT U12887 ( .A(n12315), .Y(n12757) );
  INVX1_RVT U12888 ( .A(n12315), .Y(n12758) );
  INVX1_RVT U12889 ( .A(n8313), .Y(n12759) );
  INVX1_RVT U12890 ( .A(n8313), .Y(n12760) );
  INVX1_RVT U12891 ( .A(n12326), .Y(n12761) );
  INVX1_RVT U12892 ( .A(n12324), .Y(n12762) );
  INVX1_RVT U12893 ( .A(n12325), .Y(n12763) );
  INVX1_RVT U12894 ( .A(n8165), .Y(n12764) );
  INVX1_RVT U12895 ( .A(n8165), .Y(n12765) );
  INVX1_RVT U12896 ( .A(n8262), .Y(n12766) );
  INVX1_RVT U12897 ( .A(n8262), .Y(n12767) );
  INVX1_RVT U12898 ( .A(n8209), .Y(n12768) );
  INVX1_RVT U12899 ( .A(n8209), .Y(n12769) );
  INVX1_RVT U12900 ( .A(n12313), .Y(n12770) );
  INVX1_RVT U12901 ( .A(n12350), .Y(n12771) );
  INVX1_RVT U12902 ( .A(n7357), .Y(n12772) );
  INVX1_RVT U12903 ( .A(n12348), .Y(n12773) );
  INVX1_RVT U12904 ( .A(n12348), .Y(n12774) );
  INVX1_RVT U12905 ( .A(n7482), .Y(n12775) );
  INVX1_RVT U12906 ( .A(n7482), .Y(n12776) );
  INVX1_RVT U12907 ( .A(n12359), .Y(n12777) );
  INVX1_RVT U12908 ( .A(n12357), .Y(n12778) );
  INVX1_RVT U12909 ( .A(n12358), .Y(n12779) );
  INVX1_RVT U12910 ( .A(n7334), .Y(n12780) );
  INVX1_RVT U12911 ( .A(n7334), .Y(n12781) );
  INVX1_RVT U12912 ( .A(n7431), .Y(n12782) );
  INVX1_RVT U12913 ( .A(n7431), .Y(n12783) );
  INVX1_RVT U12914 ( .A(n7378), .Y(n12784) );
  INVX1_RVT U12915 ( .A(n7378), .Y(n12785) );
  INVX1_RVT U12916 ( .A(n12346), .Y(n12786) );
  INVX1_RVT U12917 ( .A(n12383), .Y(n12787) );
  INVX1_RVT U12918 ( .A(n6518), .Y(n12788) );
  INVX1_RVT U12919 ( .A(n12381), .Y(n12789) );
  INVX1_RVT U12920 ( .A(n12381), .Y(n12790) );
  INVX1_RVT U12921 ( .A(n6643), .Y(n12791) );
  INVX1_RVT U12922 ( .A(n6643), .Y(n12792) );
  INVX1_RVT U12923 ( .A(n12392), .Y(n12793) );
  INVX1_RVT U12924 ( .A(n12390), .Y(n12794) );
  INVX1_RVT U12925 ( .A(n12391), .Y(n12795) );
  INVX1_RVT U12926 ( .A(n6495), .Y(n12796) );
  INVX1_RVT U12927 ( .A(n6495), .Y(n12797) );
  INVX1_RVT U12928 ( .A(n6592), .Y(n12798) );
  INVX1_RVT U12929 ( .A(n6592), .Y(n12799) );
  INVX1_RVT U12930 ( .A(n6539), .Y(n12800) );
  INVX1_RVT U12931 ( .A(n6539), .Y(n12801) );
  INVX1_RVT U12932 ( .A(n12379), .Y(n12802) );
  INVX1_RVT U12933 ( .A(n12647), .Y(n12803) );
  INVX1_RVT U12934 ( .A(n379), .Y(n12804) );
  INVX1_RVT U12935 ( .A(n12645), .Y(n12805) );
  INVX1_RVT U12936 ( .A(n12645), .Y(n12806) );
  INVX1_RVT U12937 ( .A(n504), .Y(n12807) );
  INVX1_RVT U12938 ( .A(n504), .Y(n12808) );
  INVX1_RVT U12939 ( .A(n12656), .Y(n12809) );
  INVX1_RVT U12940 ( .A(n12654), .Y(n12810) );
  INVX1_RVT U12941 ( .A(n12655), .Y(n12811) );
  INVX1_RVT U12942 ( .A(n356), .Y(n12812) );
  INVX1_RVT U12943 ( .A(n356), .Y(n12813) );
  INVX1_RVT U12944 ( .A(n453), .Y(n12814) );
  INVX1_RVT U12945 ( .A(n453), .Y(n12815) );
  INVX1_RVT U12946 ( .A(n400), .Y(n12816) );
  INVX1_RVT U12947 ( .A(n400), .Y(n12817) );
  INVX1_RVT U12948 ( .A(n12643), .Y(n12818) );
  INVX1_RVT U12949 ( .A(n12156), .Y(n12819) );
  INVX1_RVT U12950 ( .A(n11392), .Y(n12820) );
  INVX1_RVT U12951 ( .A(n12154), .Y(n12821) );
  INVX1_RVT U12952 ( .A(n12154), .Y(n12822) );
  INVX1_RVT U12953 ( .A(n11517), .Y(n12823) );
  INVX1_RVT U12954 ( .A(n11517), .Y(n12824) );
  INVX1_RVT U12955 ( .A(n12165), .Y(n12825) );
  INVX1_RVT U12956 ( .A(n12163), .Y(n12826) );
  INVX1_RVT U12957 ( .A(n12164), .Y(n12827) );
  INVX1_RVT U12958 ( .A(n11369), .Y(n12828) );
  INVX1_RVT U12959 ( .A(n11369), .Y(n12829) );
  INVX1_RVT U12960 ( .A(n11466), .Y(n12830) );
  INVX1_RVT U12961 ( .A(n11466), .Y(n12831) );
  INVX1_RVT U12962 ( .A(n11413), .Y(n12832) );
  INVX1_RVT U12963 ( .A(n11413), .Y(n12833) );
  INVX1_RVT U12964 ( .A(n12152), .Y(n12834) );
  INVX1_RVT U12965 ( .A(n12218), .Y(n12835) );
  INVX1_RVT U12966 ( .A(n10571), .Y(n12836) );
  INVX1_RVT U12967 ( .A(n12216), .Y(n12837) );
  INVX1_RVT U12968 ( .A(n12216), .Y(n12838) );
  INVX1_RVT U12969 ( .A(n10696), .Y(n12839) );
  INVX1_RVT U12970 ( .A(n10696), .Y(n12840) );
  INVX1_RVT U12971 ( .A(n12227), .Y(n12841) );
  INVX1_RVT U12972 ( .A(n12225), .Y(n12842) );
  INVX1_RVT U12973 ( .A(n12226), .Y(n12843) );
  INVX1_RVT U12974 ( .A(n10548), .Y(n12844) );
  INVX1_RVT U12975 ( .A(n10548), .Y(n12845) );
  INVX1_RVT U12976 ( .A(n10645), .Y(n12846) );
  INVX1_RVT U12977 ( .A(n10645), .Y(n12847) );
  INVX1_RVT U12978 ( .A(n10592), .Y(n12848) );
  INVX1_RVT U12979 ( .A(n10592), .Y(n12849) );
  INVX1_RVT U12980 ( .A(n12214), .Y(n12850) );
  INVX1_RVT U12981 ( .A(n12251), .Y(n12851) );
  INVX1_RVT U12982 ( .A(n9752), .Y(n12852) );
  INVX1_RVT U12983 ( .A(n12249), .Y(n12853) );
  INVX1_RVT U12984 ( .A(n12249), .Y(n12854) );
  INVX1_RVT U12985 ( .A(n9877), .Y(n12855) );
  INVX1_RVT U12986 ( .A(n9877), .Y(n12856) );
  INVX1_RVT U12987 ( .A(n12260), .Y(n12857) );
  INVX1_RVT U12988 ( .A(n12258), .Y(n12858) );
  INVX1_RVT U12989 ( .A(n12259), .Y(n12859) );
  INVX1_RVT U12990 ( .A(n9729), .Y(n12860) );
  INVX1_RVT U12991 ( .A(n9729), .Y(n12861) );
  INVX1_RVT U12992 ( .A(n9826), .Y(n12862) );
  INVX1_RVT U12993 ( .A(n9826), .Y(n12863) );
  INVX1_RVT U12994 ( .A(n9773), .Y(n12864) );
  INVX1_RVT U12995 ( .A(n9773), .Y(n12865) );
  INVX1_RVT U12996 ( .A(n12247), .Y(n12866) );
  INVX1_RVT U12997 ( .A(n6183), .Y(n12867) );
  INVX1_RVT U12998 ( .A(n6183), .Y(n12868) );
  INVX1_RVT U12999 ( .A(n8100), .Y(n12869) );
  INVX1_RVT U13000 ( .A(n8100), .Y(n12870) );
  INVX1_RVT U13001 ( .A(n12189), .Y(n12871) );
  INVX1_RVT U13002 ( .A(n1309), .Y(n12872) );
  INVX1_RVT U13003 ( .A(n12194), .Y(n12873) );
  INVX1_RVT U13004 ( .A(n12194), .Y(n12874) );
  INVX1_RVT U13005 ( .A(n7012), .Y(n12875) );
  INVX1_RVT U13006 ( .A(n7012), .Y(n12876) );
  INVX1_RVT U13007 ( .A(n7012), .Y(n12877) );
  INVX1_RVT U13008 ( .A(n12482), .Y(n12878) );
  INVX1_RVT U13009 ( .A(n2718), .Y(n12879) );
  INVX1_RVT U13010 ( .A(n12480), .Y(n12880) );
  INVX1_RVT U13011 ( .A(n12480), .Y(n12881) );
  INVX1_RVT U13012 ( .A(n2843), .Y(n12882) );
  INVX1_RVT U13013 ( .A(n2843), .Y(n12883) );
  INVX1_RVT U13014 ( .A(n12491), .Y(n12884) );
  INVX1_RVT U13015 ( .A(n12489), .Y(n12885) );
  INVX1_RVT U13016 ( .A(n12490), .Y(n12886) );
  INVX1_RVT U13017 ( .A(n2695), .Y(n12887) );
  INVX1_RVT U13018 ( .A(n2695), .Y(n12888) );
  INVX1_RVT U13019 ( .A(n2792), .Y(n12889) );
  INVX1_RVT U13020 ( .A(n2792), .Y(n12890) );
  INVX1_RVT U13021 ( .A(n2739), .Y(n12891) );
  INVX1_RVT U13022 ( .A(n2739), .Y(n12892) );
  INVX1_RVT U13023 ( .A(n12478), .Y(n12893) );
  INVX1_RVT U13024 ( .A(n12581), .Y(n12894) );
  INVX1_RVT U13025 ( .A(n1978), .Y(n12895) );
  INVX1_RVT U13026 ( .A(n12579), .Y(n12896) );
  INVX1_RVT U13027 ( .A(n12579), .Y(n12897) );
  INVX1_RVT U13028 ( .A(n2103), .Y(n12898) );
  INVX1_RVT U13029 ( .A(n2103), .Y(n12899) );
  INVX1_RVT U13030 ( .A(n12590), .Y(n12900) );
  INVX1_RVT U13031 ( .A(n12588), .Y(n12901) );
  INVX1_RVT U13032 ( .A(n12589), .Y(n12902) );
  INVX1_RVT U13033 ( .A(n1955), .Y(n12903) );
  INVX1_RVT U13034 ( .A(n1955), .Y(n12904) );
  INVX1_RVT U13035 ( .A(n2052), .Y(n12905) );
  INVX1_RVT U13036 ( .A(n2052), .Y(n12906) );
  INVX1_RVT U13037 ( .A(n1999), .Y(n12907) );
  INVX1_RVT U13038 ( .A(n1999), .Y(n12908) );
  INVX1_RVT U13039 ( .A(n12577), .Y(n12909) );
  INVX1_RVT U13040 ( .A(n12614), .Y(n12910) );
  INVX1_RVT U13041 ( .A(n1119), .Y(n12911) );
  INVX1_RVT U13042 ( .A(n12612), .Y(n12912) );
  INVX1_RVT U13043 ( .A(n12612), .Y(n12913) );
  INVX1_RVT U13044 ( .A(n1244), .Y(n12914) );
  INVX1_RVT U13045 ( .A(n1244), .Y(n12915) );
  INVX1_RVT U13046 ( .A(n12623), .Y(n12916) );
  INVX1_RVT U13047 ( .A(n12621), .Y(n12917) );
  INVX1_RVT U13048 ( .A(n12622), .Y(n12918) );
  INVX1_RVT U13049 ( .A(n1096), .Y(n12919) );
  INVX1_RVT U13050 ( .A(n1096), .Y(n12920) );
  INVX1_RVT U13051 ( .A(n1193), .Y(n12921) );
  INVX1_RVT U13052 ( .A(n1193), .Y(n12922) );
  INVX1_RVT U13053 ( .A(n1140), .Y(n12923) );
  INVX1_RVT U13054 ( .A(n1140), .Y(n12924) );
  INVX1_RVT U13055 ( .A(n12610), .Y(n12925) );
  INVX1_RVT U13056 ( .A(n12927), .Y(n12926) );
  INVX1_RVT U13057 ( .A(n1314), .Y(n12927) );
  INVX1_RVT U13058 ( .A(n1334), .Y(n12928) );
endmodule

