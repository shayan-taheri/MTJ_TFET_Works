module aes_16(clk, state, key, out);

    input         clk;
    input  [15:0] state, key;
    output reg [15:0] out;
				   
    reg [3:0]   p00, p01,
                p10, p11;
				
    reg [3:0]   y00, y01,
                y10, y11;
				
    reg [7:0]   k0, k1, k1x, k0_o, k1_o;
	
    wire [7:0]  k0_i, k1_i, v0, v1;

    wire [7:0]  s0,  s1,
                z0,  z1,
		g0,  g1;

    assign {s0, s1} = state ^ key;
	
    assign {k0_i, k1_i} = key;
	
    assign v0 = {k0_i[7:6] ^ 2'h1, k0_i[5:0]};
    assign v1 = v0 ^ k1_i;

    // ************* First Round *************
	
    always @ (state, key)
	
    begin
	
    {k0, k1} <= key;
	
    // First Portion
    case (s0)
    8'h00: {p00, p01} <= 8'h63;
    8'h01: {p00, p01} <= 8'h7c;
    8'h02: {p00, p01} <= 8'h77;
    8'h03: {p00, p01} <= 8'h7b;
    8'h04: {p00, p01} <= 8'hf2;
    8'h05: {p00, p01} <= 8'h6b;
    8'h06: {p00, p01} <= 8'h6f;
    8'h07: {p00, p01} <= 8'hc5;
    8'h08: {p00, p01} <= 8'h30;
    8'h09: {p00, p01} <= 8'h01;
    8'h0a: {p00, p01} <= 8'h67;
    8'h0b: {p00, p01} <= 8'h2b;
    8'h0c: {p00, p01} <= 8'hfe;
    8'h0d: {p00, p01} <= 8'hd7;
    8'h0e: {p00, p01} <= 8'hab;
    8'h0f: {p00, p01} <= 8'h76;
    8'h10: {p00, p01} <= 8'hca;
    8'h11: {p00, p01} <= 8'h82;
    8'h12: {p00, p01} <= 8'hc9;
    8'h13: {p00, p01} <= 8'h7d;
    8'h14: {p00, p01} <= 8'hfa;
    8'h15: {p00, p01} <= 8'h59;
    8'h16: {p00, p01} <= 8'h47;
    8'h17: {p00, p01} <= 8'hf0;
    8'h18: {p00, p01} <= 8'had;
    8'h19: {p00, p01} <= 8'hd4;
    8'h1a: {p00, p01} <= 8'ha2;
    8'h1b: {p00, p01} <= 8'haf;
    8'h1c: {p00, p01} <= 8'h9c;
    8'h1d: {p00, p01} <= 8'ha4;
    8'h1e: {p00, p01} <= 8'h72;
    8'h1f: {p00, p01} <= 8'hc0;
    8'h20: {p00, p01} <= 8'hb7;
    8'h21: {p00, p01} <= 8'hfd;
    8'h22: {p00, p01} <= 8'h93;
    8'h23: {p00, p01} <= 8'h26;
    8'h24: {p00, p01} <= 8'h36;
    8'h25: {p00, p01} <= 8'h3f;
    8'h26: {p00, p01} <= 8'hf7;
    8'h27: {p00, p01} <= 8'hcc;
    8'h28: {p00, p01} <= 8'h34;
    8'h29: {p00, p01} <= 8'ha5;
    8'h2a: {p00, p01} <= 8'he5;
    8'h2b: {p00, p01} <= 8'hf1;
    8'h2c: {p00, p01} <= 8'h71;
    8'h2d: {p00, p01} <= 8'hd8;
    8'h2e: {p00, p01} <= 8'h31;
    8'h2f: {p00, p01} <= 8'h15;
    8'h30: {p00, p01} <= 8'h04;
    8'h31: {p00, p01} <= 8'hc7;
    8'h32: {p00, p01} <= 8'h23;
    8'h33: {p00, p01} <= 8'hc3;
    8'h34: {p00, p01} <= 8'h18;
    8'h35: {p00, p01} <= 8'h96;
    8'h36: {p00, p01} <= 8'h05;
    8'h37: {p00, p01} <= 8'h9a;
    8'h38: {p00, p01} <= 8'h07;
    8'h39: {p00, p01} <= 8'h12;
    8'h3a: {p00, p01} <= 8'h80;
    8'h3b: {p00, p01} <= 8'he2;
    8'h3c: {p00, p01} <= 8'heb;
    8'h3d: {p00, p01} <= 8'h27;
    8'h3e: {p00, p01} <= 8'hb2;
    8'h3f: {p00, p01} <= 8'h75;
    8'h40: {p00, p01} <= 8'h09;
    8'h41: {p00, p01} <= 8'h83;
    8'h42: {p00, p01} <= 8'h2c;
    8'h43: {p00, p01} <= 8'h1a;
    8'h44: {p00, p01} <= 8'h1b;
    8'h45: {p00, p01} <= 8'h6e;
    8'h46: {p00, p01} <= 8'h5a;
    8'h47: {p00, p01} <= 8'ha0;
    8'h48: {p00, p01} <= 8'h52;
    8'h49: {p00, p01} <= 8'h3b;
    8'h4a: {p00, p01} <= 8'hd6;
    8'h4b: {p00, p01} <= 8'hb3;
    8'h4c: {p00, p01} <= 8'h29;
    8'h4d: {p00, p01} <= 8'he3;
    8'h4e: {p00, p01} <= 8'h2f;
    8'h4f: {p00, p01} <= 8'h84;
    8'h50: {p00, p01} <= 8'h53;
    8'h51: {p00, p01} <= 8'hd1;
    8'h52: {p00, p01} <= 8'h00;
    8'h53: {p00, p01} <= 8'hed;
    8'h54: {p00, p01} <= 8'h20;
    8'h55: {p00, p01} <= 8'hfc;
    8'h56: {p00, p01} <= 8'hb1;
    8'h57: {p00, p01} <= 8'h5b;
    8'h58: {p00, p01} <= 8'h6a;
    8'h59: {p00, p01} <= 8'hcb;
    8'h5a: {p00, p01} <= 8'hbe;
    8'h5b: {p00, p01} <= 8'h39;
    8'h5c: {p00, p01} <= 8'h4a;
    8'h5d: {p00, p01} <= 8'h4c;
    8'h5e: {p00, p01} <= 8'h58;
    8'h5f: {p00, p01} <= 8'hcf;
    8'h60: {p00, p01} <= 8'hd0;
    8'h61: {p00, p01} <= 8'hef;
    8'h62: {p00, p01} <= 8'haa;
    8'h63: {p00, p01} <= 8'hfb;
    8'h64: {p00, p01} <= 8'h43;
    8'h65: {p00, p01} <= 8'h4d;
    8'h66: {p00, p01} <= 8'h33;
    8'h67: {p00, p01} <= 8'h85;
    8'h68: {p00, p01} <= 8'h45;
    8'h69: {p00, p01} <= 8'hf9;
    8'h6a: {p00, p01} <= 8'h02;
    8'h6b: {p00, p01} <= 8'h7f;
    8'h6c: {p00, p01} <= 8'h50;
    8'h6d: {p00, p01} <= 8'h3c;
    8'h6e: {p00, p01} <= 8'h9f;
    8'h6f: {p00, p01} <= 8'ha8;
    8'h70: {p00, p01} <= 8'h51;
    8'h71: {p00, p01} <= 8'ha3;
    8'h72: {p00, p01} <= 8'h40;
    8'h73: {p00, p01} <= 8'h8f;
    8'h74: {p00, p01} <= 8'h92;
    8'h75: {p00, p01} <= 8'h9d;
    8'h76: {p00, p01} <= 8'h38;
    8'h77: {p00, p01} <= 8'hf5;
    8'h78: {p00, p01} <= 8'hbc;
    8'h79: {p00, p01} <= 8'hb6;
    8'h7a: {p00, p01} <= 8'hda;
    8'h7b: {p00, p01} <= 8'h21;
    8'h7c: {p00, p01} <= 8'h10;
    8'h7d: {p00, p01} <= 8'hff;
    8'h7e: {p00, p01} <= 8'hf3;
    8'h7f: {p00, p01} <= 8'hd2;
    8'h80: {p00, p01} <= 8'hcd;
    8'h81: {p00, p01} <= 8'h0c;
    8'h82: {p00, p01} <= 8'h13;
    8'h83: {p00, p01} <= 8'hec;
    8'h84: {p00, p01} <= 8'h5f;
    8'h85: {p00, p01} <= 8'h97;
    8'h86: {p00, p01} <= 8'h44;
    8'h87: {p00, p01} <= 8'h17;
    8'h88: {p00, p01} <= 8'hc4;
    8'h89: {p00, p01} <= 8'ha7;
    8'h8a: {p00, p01} <= 8'h7e;
    8'h8b: {p00, p01} <= 8'h3d;
    8'h8c: {p00, p01} <= 8'h64;
    8'h8d: {p00, p01} <= 8'h5d;
    8'h8e: {p00, p01} <= 8'h19;
    8'h8f: {p00, p01} <= 8'h73;
    8'h90: {p00, p01} <= 8'h60;
    8'h91: {p00, p01} <= 8'h81;
    8'h92: {p00, p01} <= 8'h4f;
    8'h93: {p00, p01} <= 8'hdc;
    8'h94: {p00, p01} <= 8'h22;
    8'h95: {p00, p01} <= 8'h2a;
    8'h96: {p00, p01} <= 8'h90;
    8'h97: {p00, p01} <= 8'h88;
    8'h98: {p00, p01} <= 8'h46;
    8'h99: {p00, p01} <= 8'hee;
    8'h9a: {p00, p01} <= 8'hb8;
    8'h9b: {p00, p01} <= 8'h14;
    8'h9c: {p00, p01} <= 8'hde;
    8'h9d: {p00, p01} <= 8'h5e;
    8'h9e: {p00, p01} <= 8'h0b;
    8'h9f: {p00, p01} <= 8'hdb;
    8'ha0: {p00, p01} <= 8'he0;
    8'ha1: {p00, p01} <= 8'h32;
    8'ha2: {p00, p01} <= 8'h3a;
    8'ha3: {p00, p01} <= 8'h0a;
    8'ha4: {p00, p01} <= 8'h49;
    8'ha5: {p00, p01} <= 8'h06;
    8'ha6: {p00, p01} <= 8'h24;
    8'ha7: {p00, p01} <= 8'h5c;
    8'ha8: {p00, p01} <= 8'hc2;
    8'ha9: {p00, p01} <= 8'hd3;
    8'haa: {p00, p01} <= 8'hac;
    8'hab: {p00, p01} <= 8'h62;
    8'hac: {p00, p01} <= 8'h91;
    8'had: {p00, p01} <= 8'h95;
    8'hae: {p00, p01} <= 8'he4;
    8'haf: {p00, p01} <= 8'h79;
    8'hb0: {p00, p01} <= 8'he7;
    8'hb1: {p00, p01} <= 8'hc8;
    8'hb2: {p00, p01} <= 8'h37;
    8'hb3: {p00, p01} <= 8'h6d;
    8'hb4: {p00, p01} <= 8'h8d;
    8'hb5: {p00, p01} <= 8'hd5;
    8'hb6: {p00, p01} <= 8'h4e;
    8'hb7: {p00, p01} <= 8'ha9;
    8'hb8: {p00, p01} <= 8'h6c;
    8'hb9: {p00, p01} <= 8'h56;
    8'hba: {p00, p01} <= 8'hf4;
    8'hbb: {p00, p01} <= 8'hea;
    8'hbc: {p00, p01} <= 8'h65;
    8'hbd: {p00, p01} <= 8'h7a;
    8'hbe: {p00, p01} <= 8'hae;
    8'hbf: {p00, p01} <= 8'h08;
    8'hc0: {p00, p01} <= 8'hba;
    8'hc1: {p00, p01} <= 8'h78;
    8'hc2: {p00, p01} <= 8'h25;
    8'hc3: {p00, p01} <= 8'h2e;
    8'hc4: {p00, p01} <= 8'h1c;
    8'hc5: {p00, p01} <= 8'ha6;
    8'hc6: {p00, p01} <= 8'hb4;
    8'hc7: {p00, p01} <= 8'hc6;
    8'hc8: {p00, p01} <= 8'he8;
    8'hc9: {p00, p01} <= 8'hdd;
    8'hca: {p00, p01} <= 8'h74;
    8'hcb: {p00, p01} <= 8'h1f;
    8'hcc: {p00, p01} <= 8'h4b;
    8'hcd: {p00, p01} <= 8'hbd;
    8'hce: {p00, p01} <= 8'h8b;
    8'hcf: {p00, p01} <= 8'h8a;
    8'hd0: {p00, p01} <= 8'h70;
    8'hd1: {p00, p01} <= 8'h3e;
    8'hd2: {p00, p01} <= 8'hb5;
    8'hd3: {p00, p01} <= 8'h66;
    8'hd4: {p00, p01} <= 8'h48;
    8'hd5: {p00, p01} <= 8'h03;
    8'hd6: {p00, p01} <= 8'hf6;
    8'hd7: {p00, p01} <= 8'h0e;
    8'hd8: {p00, p01} <= 8'h61;
    8'hd9: {p00, p01} <= 8'h35;
    8'hda: {p00, p01} <= 8'h57;
    8'hdb: {p00, p01} <= 8'hb9;
    8'hdc: {p00, p01} <= 8'h86;
    8'hdd: {p00, p01} <= 8'hc1;
    8'hde: {p00, p01} <= 8'h1d;
    8'hdf: {p00, p01} <= 8'h9e;
    8'he0: {p00, p01} <= 8'he1;
    8'he1: {p00, p01} <= 8'hf8;
    8'he2: {p00, p01} <= 8'h98;
    8'he3: {p00, p01} <= 8'h11;
    8'he4: {p00, p01} <= 8'h69;
    8'he5: {p00, p01} <= 8'hd9;
    8'he6: {p00, p01} <= 8'h8e;
    8'he7: {p00, p01} <= 8'h94;
    8'he8: {p00, p01} <= 8'h9b;
    8'he9: {p00, p01} <= 8'h1e;
    8'hea: {p00, p01} <= 8'h87;
    8'heb: {p00, p01} <= 8'he9;
    8'hec: {p00, p01} <= 8'hce;
    8'hed: {p00, p01} <= 8'h55;
    8'hee: {p00, p01} <= 8'h28;
    8'hef: {p00, p01} <= 8'hdf;
    8'hf0: {p00, p01} <= 8'h8c;
    8'hf1: {p00, p01} <= 8'ha1;
    8'hf2: {p00, p01} <= 8'h89;
    8'hf3: {p00, p01} <= 8'h0d;
    8'hf4: {p00, p01} <= 8'hbf;
    8'hf5: {p00, p01} <= 8'he6;
    8'hf6: {p00, p01} <= 8'h42;
    8'hf7: {p00, p01} <= 8'h68;
    8'hf8: {p00, p01} <= 8'h41;
    8'hf9: {p00, p01} <= 8'h99;
    8'hfa: {p00, p01} <= 8'h2d;
    8'hfb: {p00, p01} <= 8'h0f;
    8'hfc: {p00, p01} <= 8'hb0;
    8'hfd: {p00, p01} <= 8'h54;
    8'hfe: {p00, p01} <= 8'hbb;
    8'hff: {p00, p01} <= 8'h16;
    endcase
	
	
	
	
    // Second Portion
    case (s1)
    8'h00: {p10, p11} <= 8'h63;
    8'h01: {p10, p11} <= 8'h7c;
    8'h02: {p10, p11} <= 8'h77;
    8'h03: {p10, p11} <= 8'h7b;
    8'h04: {p10, p11} <= 8'hf2;
    8'h05: {p10, p11} <= 8'h6b;
    8'h06: {p10, p11} <= 8'h6f;
    8'h07: {p10, p11} <= 8'hc5;
    8'h08: {p10, p11} <= 8'h30;
    8'h09: {p10, p11} <= 8'h01;
    8'h0a: {p10, p11} <= 8'h67;
    8'h0b: {p10, p11} <= 8'h2b;
    8'h0c: {p10, p11} <= 8'hfe;
    8'h0d: {p10, p11} <= 8'hd7;
    8'h0e: {p10, p11} <= 8'hab;
    8'h0f: {p10, p11} <= 8'h76;
    8'h10: {p10, p11} <= 8'hca;
    8'h11: {p10, p11} <= 8'h82;
    8'h12: {p10, p11} <= 8'hc9;
    8'h13: {p10, p11} <= 8'h7d;
    8'h14: {p10, p11} <= 8'hfa;
    8'h15: {p10, p11} <= 8'h59;
    8'h16: {p10, p11} <= 8'h47;
    8'h17: {p10, p11} <= 8'hf0;
    8'h18: {p10, p11} <= 8'had;
    8'h19: {p10, p11} <= 8'hd4;
    8'h1a: {p10, p11} <= 8'ha2;
    8'h1b: {p10, p11} <= 8'haf;
    8'h1c: {p10, p11} <= 8'h9c;
    8'h1d: {p10, p11} <= 8'ha4;
    8'h1e: {p10, p11} <= 8'h72;
    8'h1f: {p10, p11} <= 8'hc0;
    8'h20: {p10, p11} <= 8'hb7;
    8'h21: {p10, p11} <= 8'hfd;
    8'h22: {p10, p11} <= 8'h93;
    8'h23: {p10, p11} <= 8'h26;
    8'h24: {p10, p11} <= 8'h36;
    8'h25: {p10, p11} <= 8'h3f;
    8'h26: {p10, p11} <= 8'hf7;
    8'h27: {p10, p11} <= 8'hcc;
    8'h28: {p10, p11} <= 8'h34;
    8'h29: {p10, p11} <= 8'ha5;
    8'h2a: {p10, p11} <= 8'he5;
    8'h2b: {p10, p11} <= 8'hf1;
    8'h2c: {p10, p11} <= 8'h71;
    8'h2d: {p10, p11} <= 8'hd8;
    8'h2e: {p10, p11} <= 8'h31;
    8'h2f: {p10, p11} <= 8'h15;
    8'h30: {p10, p11} <= 8'h04;
    8'h31: {p10, p11} <= 8'hc7;
    8'h32: {p10, p11} <= 8'h23;
    8'h33: {p10, p11} <= 8'hc3;
    8'h34: {p10, p11} <= 8'h18;
    8'h35: {p10, p11} <= 8'h96;
    8'h36: {p10, p11} <= 8'h05;
    8'h37: {p10, p11} <= 8'h9a;
    8'h38: {p10, p11} <= 8'h07;
    8'h39: {p10, p11} <= 8'h12;
    8'h3a: {p10, p11} <= 8'h80;
    8'h3b: {p10, p11} <= 8'he2;
    8'h3c: {p10, p11} <= 8'heb;
    8'h3d: {p10, p11} <= 8'h27;
    8'h3e: {p10, p11} <= 8'hb2;
    8'h3f: {p10, p11} <= 8'h75;
    8'h40: {p10, p11} <= 8'h09;
    8'h41: {p10, p11} <= 8'h83;
    8'h42: {p10, p11} <= 8'h2c;
    8'h43: {p10, p11} <= 8'h1a;
    8'h44: {p10, p11} <= 8'h1b;
    8'h45: {p10, p11} <= 8'h6e;
    8'h46: {p10, p11} <= 8'h5a;
    8'h47: {p10, p11} <= 8'ha0;
    8'h48: {p10, p11} <= 8'h52;
    8'h49: {p10, p11} <= 8'h3b;
    8'h4a: {p10, p11} <= 8'hd6;
    8'h4b: {p10, p11} <= 8'hb3;
    8'h4c: {p10, p11} <= 8'h29;
    8'h4d: {p10, p11} <= 8'he3;
    8'h4e: {p10, p11} <= 8'h2f;
    8'h4f: {p10, p11} <= 8'h84;
    8'h50: {p10, p11} <= 8'h53;
    8'h51: {p10, p11} <= 8'hd1;
    8'h52: {p10, p11} <= 8'h00;
    8'h53: {p10, p11} <= 8'hed;
    8'h54: {p10, p11} <= 8'h20;
    8'h55: {p10, p11} <= 8'hfc;
    8'h56: {p10, p11} <= 8'hb1;
    8'h57: {p10, p11} <= 8'h5b;
    8'h58: {p10, p11} <= 8'h6a;
    8'h59: {p10, p11} <= 8'hcb;
    8'h5a: {p10, p11} <= 8'hbe;
    8'h5b: {p10, p11} <= 8'h39;
    8'h5c: {p10, p11} <= 8'h4a;
    8'h5d: {p10, p11} <= 8'h4c;
    8'h5e: {p10, p11} <= 8'h58;
    8'h5f: {p10, p11} <= 8'hcf;
    8'h60: {p10, p11} <= 8'hd0;
    8'h61: {p10, p11} <= 8'hef;
    8'h62: {p10, p11} <= 8'haa;
    8'h63: {p10, p11} <= 8'hfb;
    8'h64: {p10, p11} <= 8'h43;
    8'h65: {p10, p11} <= 8'h4d;
    8'h66: {p10, p11} <= 8'h33;
    8'h67: {p10, p11} <= 8'h85;
    8'h68: {p10, p11} <= 8'h45;
    8'h69: {p10, p11} <= 8'hf9;
    8'h6a: {p10, p11} <= 8'h02;
    8'h6b: {p10, p11} <= 8'h7f;
    8'h6c: {p10, p11} <= 8'h50;
    8'h6d: {p10, p11} <= 8'h3c;
    8'h6e: {p10, p11} <= 8'h9f;
    8'h6f: {p10, p11} <= 8'ha8;
    8'h70: {p10, p11} <= 8'h51;
    8'h71: {p10, p11} <= 8'ha3;
    8'h72: {p10, p11} <= 8'h40;
    8'h73: {p10, p11} <= 8'h8f;
    8'h74: {p10, p11} <= 8'h92;
    8'h75: {p10, p11} <= 8'h9d;
    8'h76: {p10, p11} <= 8'h38;
    8'h77: {p10, p11} <= 8'hf5;
    8'h78: {p10, p11} <= 8'hbc;
    8'h79: {p10, p11} <= 8'hb6;
    8'h7a: {p10, p11} <= 8'hda;
    8'h7b: {p10, p11} <= 8'h21;
    8'h7c: {p10, p11} <= 8'h10;
    8'h7d: {p10, p11} <= 8'hff;
    8'h7e: {p10, p11} <= 8'hf3;
    8'h7f: {p10, p11} <= 8'hd2;
    8'h80: {p10, p11} <= 8'hcd;
    8'h81: {p10, p11} <= 8'h0c;
    8'h82: {p10, p11} <= 8'h13;
    8'h83: {p10, p11} <= 8'hec;
    8'h84: {p10, p11} <= 8'h5f;
    8'h85: {p10, p11} <= 8'h97;
    8'h86: {p10, p11} <= 8'h44;
    8'h87: {p10, p11} <= 8'h17;
    8'h88: {p10, p11} <= 8'hc4;
    8'h89: {p10, p11} <= 8'ha7;
    8'h8a: {p10, p11} <= 8'h7e;
    8'h8b: {p10, p11} <= 8'h3d;
    8'h8c: {p10, p11} <= 8'h64;
    8'h8d: {p10, p11} <= 8'h5d;
    8'h8e: {p10, p11} <= 8'h19;
    8'h8f: {p10, p11} <= 8'h73;
    8'h90: {p10, p11} <= 8'h60;
    8'h91: {p10, p11} <= 8'h81;
    8'h92: {p10, p11} <= 8'h4f;
    8'h93: {p10, p11} <= 8'hdc;
    8'h94: {p10, p11} <= 8'h22;
    8'h95: {p10, p11} <= 8'h2a;
    8'h96: {p10, p11} <= 8'h90;
    8'h97: {p10, p11} <= 8'h88;
    8'h98: {p10, p11} <= 8'h46;
    8'h99: {p10, p11} <= 8'hee;
    8'h9a: {p10, p11} <= 8'hb8;
    8'h9b: {p10, p11} <= 8'h14;
    8'h9c: {p10, p11} <= 8'hde;
    8'h9d: {p10, p11} <= 8'h5e;
    8'h9e: {p10, p11} <= 8'h0b;
    8'h9f: {p10, p11} <= 8'hdb;
    8'ha0: {p10, p11} <= 8'he0;
    8'ha1: {p10, p11} <= 8'h32;
    8'ha2: {p10, p11} <= 8'h3a;
    8'ha3: {p10, p11} <= 8'h0a;
    8'ha4: {p10, p11} <= 8'h49;
    8'ha5: {p10, p11} <= 8'h06;
    8'ha6: {p10, p11} <= 8'h24;
    8'ha7: {p10, p11} <= 8'h5c;
    8'ha8: {p10, p11} <= 8'hc2;
    8'ha9: {p10, p11} <= 8'hd3;
    8'haa: {p10, p11} <= 8'hac;
    8'hab: {p10, p11} <= 8'h62;
    8'hac: {p10, p11} <= 8'h91;
    8'had: {p10, p11} <= 8'h95;
    8'hae: {p10, p11} <= 8'he4;
    8'haf: {p10, p11} <= 8'h79;
    8'hb0: {p10, p11} <= 8'he7;
    8'hb1: {p10, p11} <= 8'hc8;
    8'hb2: {p10, p11} <= 8'h37;
    8'hb3: {p10, p11} <= 8'h6d;
    8'hb4: {p10, p11} <= 8'h8d;
    8'hb5: {p10, p11} <= 8'hd5;
    8'hb6: {p10, p11} <= 8'h4e;
    8'hb7: {p10, p11} <= 8'ha9;
    8'hb8: {p10, p11} <= 8'h6c;
    8'hb9: {p10, p11} <= 8'h56;
    8'hba: {p10, p11} <= 8'hf4;
    8'hbb: {p10, p11} <= 8'hea;
    8'hbc: {p10, p11} <= 8'h65;
    8'hbd: {p10, p11} <= 8'h7a;
    8'hbe: {p10, p11} <= 8'hae;
    8'hbf: {p10, p11} <= 8'h08;
    8'hc0: {p10, p11} <= 8'hba;
    8'hc1: {p10, p11} <= 8'h78;
    8'hc2: {p10, p11} <= 8'h25;
    8'hc3: {p10, p11} <= 8'h2e;
    8'hc4: {p10, p11} <= 8'h1c;
    8'hc5: {p10, p11} <= 8'ha6;
    8'hc6: {p10, p11} <= 8'hb4;
    8'hc7: {p10, p11} <= 8'hc6;
    8'hc8: {p10, p11} <= 8'he8;
    8'hc9: {p10, p11} <= 8'hdd;
    8'hca: {p10, p11} <= 8'h74;
    8'hcb: {p10, p11} <= 8'h1f;
    8'hcc: {p10, p11} <= 8'h4b;
    8'hcd: {p10, p11} <= 8'hbd;
    8'hce: {p10, p11} <= 8'h8b;
    8'hcf: {p10, p11} <= 8'h8a;
    8'hd0: {p10, p11} <= 8'h70;
    8'hd1: {p10, p11} <= 8'h3e;
    8'hd2: {p10, p11} <= 8'hb5;
    8'hd3: {p10, p11} <= 8'h66;
    8'hd4: {p10, p11} <= 8'h48;
    8'hd5: {p10, p11} <= 8'h03;
    8'hd6: {p10, p11} <= 8'hf6;
    8'hd7: {p10, p11} <= 8'h0e;
    8'hd8: {p10, p11} <= 8'h61;
    8'hd9: {p10, p11} <= 8'h35;
    8'hda: {p10, p11} <= 8'h57;
    8'hdb: {p10, p11} <= 8'hb9;
    8'hdc: {p10, p11} <= 8'h86;
    8'hdd: {p10, p11} <= 8'hc1;
    8'hde: {p10, p11} <= 8'h1d;
    8'hdf: {p10, p11} <= 8'h9e;
    8'he0: {p10, p11} <= 8'he1;
    8'he1: {p10, p11} <= 8'hf8;
    8'he2: {p10, p11} <= 8'h98;
    8'he3: {p10, p11} <= 8'h11;
    8'he4: {p10, p11} <= 8'h69;
    8'he5: {p10, p11} <= 8'hd9;
    8'he6: {p10, p11} <= 8'h8e;
    8'he7: {p10, p11} <= 8'h94;
    8'he8: {p10, p11} <= 8'h9b;
    8'he9: {p10, p11} <= 8'h1e;
    8'hea: {p10, p11} <= 8'h87;
    8'heb: {p10, p11} <= 8'he9;
    8'hec: {p10, p11} <= 8'hce;
    8'hed: {p10, p11} <= 8'h55;
    8'hee: {p10, p11} <= 8'h28;
    8'hef: {p10, p11} <= 8'hdf;
    8'hf0: {p10, p11} <= 8'h8c;
    8'hf1: {p10, p11} <= 8'ha1;
    8'hf2: {p10, p11} <= 8'h89;
    8'hf3: {p10, p11} <= 8'h0d;
    8'hf4: {p10, p11} <= 8'hbf;
    8'hf5: {p10, p11} <= 8'he6;
    8'hf6: {p10, p11} <= 8'h42;
    8'hf7: {p10, p11} <= 8'h68;
    8'hf8: {p10, p11} <= 8'h41;
    8'hf9: {p10, p11} <= 8'h99;
    8'hfa: {p10, p11} <= 8'h2d;
    8'hfb: {p10, p11} <= 8'h0f;
    8'hfc: {p10, p11} <= 8'hb0;
    8'hfd: {p10, p11} <= 8'h54;
    8'hfe: {p10, p11} <= 8'hbb;
    8'hff: {p10, p11} <= 8'h16;
    endcase
	
    case (k1_i)
    8'h00: k1x <= 8'h63;
    8'h01: k1x <= 8'h7c;
    8'h02: k1x <= 8'h77;
    8'h03: k1x <= 8'h7b;
    8'h04: k1x <= 8'hf2;
    8'h05: k1x <= 8'h6b;
    8'h06: k1x <= 8'h6f;
    8'h07: k1x <= 8'hc5;
    8'h08: k1x <= 8'h30;
    8'h09: k1x <= 8'h01;
    8'h0a: k1x <= 8'h67;
    8'h0b: k1x <= 8'h2b;
    8'h0c: k1x <= 8'hfe;
    8'h0d: k1x <= 8'hd7;
    8'h0e: k1x <= 8'hab;
    8'h0f: k1x <= 8'h76;
    8'h10: k1x <= 8'hca;
    8'h11: k1x <= 8'h82;
    8'h12: k1x <= 8'hc9;
    8'h13: k1x <= 8'h7d;
    8'h14: k1x <= 8'hfa;
    8'h15: k1x <= 8'h59;
    8'h16: k1x <= 8'h47;
    8'h17: k1x <= 8'hf0;
    8'h18: k1x <= 8'had;
    8'h19: k1x <= 8'hd4;
    8'h1a: k1x <= 8'ha2;
    8'h1b: k1x <= 8'haf;
    8'h1c: k1x <= 8'h9c;
    8'h1d: k1x <= 8'ha4;
    8'h1e: k1x <= 8'h72;
    8'h1f: k1x <= 8'hc0;
    8'h20: k1x <= 8'hb7;
    8'h21: k1x <= 8'hfd;
    8'h22: k1x <= 8'h93;
    8'h23: k1x <= 8'h26;
    8'h24: k1x <= 8'h36;
    8'h25: k1x <= 8'h3f;
    8'h26: k1x <= 8'hf7;
    8'h27: k1x <= 8'hcc;
    8'h28: k1x <= 8'h34;
    8'h29: k1x <= 8'ha5;
    8'h2a: k1x <= 8'he5;
    8'h2b: k1x <= 8'hf1;
    8'h2c: k1x <= 8'h71;
    8'h2d: k1x <= 8'hd8;
    8'h2e: k1x <= 8'h31;
    8'h2f: k1x <= 8'h15;
    8'h30: k1x <= 8'h04;
    8'h31: k1x <= 8'hc7;
    8'h32: k1x <= 8'h23;
    8'h33: k1x <= 8'hc3;
    8'h34: k1x <= 8'h18;
    8'h35: k1x <= 8'h96;
    8'h36: k1x <= 8'h05;
    8'h37: k1x <= 8'h9a;
    8'h38: k1x <= 8'h07;
    8'h39: k1x <= 8'h12;
    8'h3a: k1x <= 8'h80;
    8'h3b: k1x <= 8'he2;
    8'h3c: k1x <= 8'heb;
    8'h3d: k1x <= 8'h27;
    8'h3e: k1x <= 8'hb2;
    8'h3f: k1x <= 8'h75;
    8'h40: k1x <= 8'h09;
    8'h41: k1x <= 8'h83;
    8'h42: k1x <= 8'h2c;
    8'h43: k1x <= 8'h1a;
    8'h44: k1x <= 8'h1b;
    8'h45: k1x <= 8'h6e;
    8'h46: k1x <= 8'h5a;
    8'h47: k1x <= 8'ha0;
    8'h48: k1x <= 8'h52;
    8'h49: k1x <= 8'h3b;
    8'h4a: k1x <= 8'hd6;
    8'h4b: k1x <= 8'hb3;
    8'h4c: k1x <= 8'h29;
    8'h4d: k1x <= 8'he3;
    8'h4e: k1x <= 8'h2f;
    8'h4f: k1x <= 8'h84;
    8'h50: k1x <= 8'h53;
    8'h51: k1x <= 8'hd1;
    8'h52: k1x <= 8'h00;
    8'h53: k1x <= 8'hed;
    8'h54: k1x <= 8'h20;
    8'h55: k1x <= 8'hfc;
    8'h56: k1x <= 8'hb1;
    8'h57: k1x <= 8'h5b;
    8'h58: k1x <= 8'h6a;
    8'h59: k1x <= 8'hcb;
    8'h5a: k1x <= 8'hbe;
    8'h5b: k1x <= 8'h39;
    8'h5c: k1x <= 8'h4a;
    8'h5d: k1x <= 8'h4c;
    8'h5e: k1x <= 8'h58;
    8'h5f: k1x <= 8'hcf;
    8'h60: k1x <= 8'hd0;
    8'h61: k1x <= 8'hef;
    8'h62: k1x <= 8'haa;
    8'h63: k1x <= 8'hfb;
    8'h64: k1x <= 8'h43;
    8'h65: k1x <= 8'h4d;
    8'h66: k1x <= 8'h33;
    8'h67: k1x <= 8'h85;
    8'h68: k1x <= 8'h45;
    8'h69: k1x <= 8'hf9;
    8'h6a: k1x <= 8'h02;
    8'h6b: k1x <= 8'h7f;
    8'h6c: k1x <= 8'h50;
    8'h6d: k1x <= 8'h3c;
    8'h6e: k1x <= 8'h9f;
    8'h6f: k1x <= 8'ha8;
    8'h70: k1x <= 8'h51;
    8'h71: k1x <= 8'ha3;
    8'h72: k1x <= 8'h40;
    8'h73: k1x <= 8'h8f;
    8'h74: k1x <= 8'h92;
    8'h75: k1x <= 8'h9d;
    8'h76: k1x <= 8'h38;
    8'h77: k1x <= 8'hf5;
    8'h78: k1x <= 8'hbc;
    8'h79: k1x <= 8'hb6;
    8'h7a: k1x <= 8'hda;
    8'h7b: k1x <= 8'h21;
    8'h7c: k1x <= 8'h10;
    8'h7d: k1x <= 8'hff;
    8'h7e: k1x <= 8'hf3;
    8'h7f: k1x <= 8'hd2;
    8'h80: k1x <= 8'hcd;
    8'h81: k1x <= 8'h0c;
    8'h82: k1x <= 8'h13;
    8'h83: k1x <= 8'hec;
    8'h84: k1x <= 8'h5f;
    8'h85: k1x <= 8'h97;
    8'h86: k1x <= 8'h44;
    8'h87: k1x <= 8'h17;
    8'h88: k1x <= 8'hc4;
    8'h89: k1x <= 8'ha7;
    8'h8a: k1x <= 8'h7e;
    8'h8b: k1x <= 8'h3d;
    8'h8c: k1x <= 8'h64;
    8'h8d: k1x <= 8'h5d;
    8'h8e: k1x <= 8'h19;
    8'h8f: k1x <= 8'h73;
    8'h90: k1x <= 8'h60;
    8'h91: k1x <= 8'h81;
    8'h92: k1x <= 8'h4f;
    8'h93: k1x <= 8'hdc;
    8'h94: k1x <= 8'h22;
    8'h95: k1x <= 8'h2a;
    8'h96: k1x <= 8'h90;
    8'h97: k1x <= 8'h88;
    8'h98: k1x <= 8'h46;
    8'h99: k1x <= 8'hee;
    8'h9a: k1x <= 8'hb8;
    8'h9b: k1x <= 8'h14;
    8'h9c: k1x <= 8'hde;
    8'h9d: k1x <= 8'h5e;
    8'h9e: k1x <= 8'h0b;
    8'h9f: k1x <= 8'hdb;
    8'ha0: k1x <= 8'he0;
    8'ha1: k1x <= 8'h32;
    8'ha2: k1x <= 8'h3a;
    8'ha3: k1x <= 8'h0a;
    8'ha4: k1x <= 8'h49;
    8'ha5: k1x <= 8'h06;
    8'ha6: k1x <= 8'h24;
    8'ha7: k1x <= 8'h5c;
    8'ha8: k1x <= 8'hc2;
    8'ha9: k1x <= 8'hd3;
    8'haa: k1x <= 8'hac;
    8'hab: k1x <= 8'h62;
    8'hac: k1x <= 8'h91;
    8'had: k1x <= 8'h95;
    8'hae: k1x <= 8'he4;
    8'haf: k1x <= 8'h79;
    8'hb0: k1x <= 8'he7;
    8'hb1: k1x <= 8'hc8;
    8'hb2: k1x <= 8'h37;
    8'hb3: k1x <= 8'h6d;
    8'hb4: k1x <= 8'h8d;
    8'hb5: k1x <= 8'hd5;
    8'hb6: k1x <= 8'h4e;
    8'hb7: k1x <= 8'ha9;
    8'hb8: k1x <= 8'h6c;
    8'hb9: k1x <= 8'h56;
    8'hba: k1x <= 8'hf4;
    8'hbb: k1x <= 8'hea;
    8'hbc: k1x <= 8'h65;
    8'hbd: k1x <= 8'h7a;
    8'hbe: k1x <= 8'hae;
    8'hbf: k1x <= 8'h08;
    8'hc0: k1x <= 8'hba;
    8'hc1: k1x <= 8'h78;
    8'hc2: k1x <= 8'h25;
    8'hc3: k1x <= 8'h2e;
    8'hc4: k1x <= 8'h1c;
    8'hc5: k1x <= 8'ha6;
    8'hc6: k1x <= 8'hb4;
    8'hc7: k1x <= 8'hc6;
    8'hc8: k1x <= 8'he8;
    8'hc9: k1x <= 8'hdd;
    8'hca: k1x <= 8'h74;
    8'hcb: k1x <= 8'h1f;
    8'hcc: k1x <= 8'h4b;
    8'hcd: k1x <= 8'hbd;
    8'hce: k1x <= 8'h8b;
    8'hcf: k1x <= 8'h8a;
    8'hd0: k1x <= 8'h70;
    8'hd1: k1x <= 8'h3e;
    8'hd2: k1x <= 8'hb5;
    8'hd3: k1x <= 8'h66;
    8'hd4: k1x <= 8'h48;
    8'hd5: k1x <= 8'h03;
    8'hd6: k1x <= 8'hf6;
    8'hd7: k1x <= 8'h0e;
    8'hd8: k1x <= 8'h61;
    8'hd9: k1x <= 8'h35;
    8'hda: k1x <= 8'h57;
    8'hdb: k1x <= 8'hb9;
    8'hdc: k1x <= 8'h86;
    8'hdd: k1x <= 8'hc1;
    8'hde: k1x <= 8'h1d;
    8'hdf: k1x <= 8'h9e;
    8'he0: k1x <= 8'he1;
    8'he1: k1x <= 8'hf8;
    8'he2: k1x <= 8'h98;
    8'he3: k1x <= 8'h11;
    8'he4: k1x <= 8'h69;
    8'he5: k1x <= 8'hd9;
    8'he6: k1x <= 8'h8e;
    8'he7: k1x <= 8'h94;
    8'he8: k1x <= 8'h9b;
    8'he9: k1x <= 8'h1e;
    8'hea: k1x <= 8'h87;
    8'heb: k1x <= 8'he9;
    8'hec: k1x <= 8'hce;
    8'hed: k1x <= 8'h55;
    8'hee: k1x <= 8'h28;
    8'hef: k1x <= 8'hdf;
    8'hf0: k1x <= 8'h8c;
    8'hf1: k1x <= 8'ha1;
    8'hf2: k1x <= 8'h89;
    8'hf3: k1x <= 8'h0d;
    8'hf4: k1x <= 8'hbf;
    8'hf5: k1x <= 8'he6;
    8'hf6: k1x <= 8'h42;
    8'hf7: k1x <= 8'h68;
    8'hf8: k1x <= 8'h41;
    8'hf9: k1x <= 8'h99;
    8'hfa: k1x <= 8'h2d;
    8'hfb: k1x <= 8'h0f;
    8'hfc: k1x <= 8'hb0;
    8'hfd: k1x <= 8'h54;
    8'hfe: k1x <= 8'hbb;
    8'hff: k1x <= 8'h16;
    endcase
	
    end

    assign z0 = {p00, p11} ^ k0;
    assign z1 = {p10, p01} ^ k1;
	
	
    // ***************************************

    // ************* Second Round *************
	
    always @ (z0, z1, k1x)
	
    begin
	
    k0_o <= v0 ^ k1x;
    k1_o <= v1 ^ k1x;
	
    case (z0)
    8'h00: {y00, y01} <= 8'h63;
    8'h01: {y00, y01} <= 8'h7c;
    8'h02: {y00, y01} <= 8'h77;
    8'h03: {y00, y01} <= 8'h7b;
    8'h04: {y00, y01} <= 8'hf2;
    8'h05: {y00, y01} <= 8'h6b;
    8'h06: {y00, y01} <= 8'h6f;
    8'h07: {y00, y01} <= 8'hc5;
    8'h08: {y00, y01} <= 8'h30;
    8'h09: {y00, y01} <= 8'h01;
    8'h0a: {y00, y01} <= 8'h67;
    8'h0b: {y00, y01} <= 8'h2b;
    8'h0c: {y00, y01} <= 8'hfe;
    8'h0d: {y00, y01} <= 8'hd7;
    8'h0e: {y00, y01} <= 8'hab;
    8'h0f: {y00, y01} <= 8'h76;
    8'h10: {y00, y01} <= 8'hca;
    8'h11: {y00, y01} <= 8'h82;
    8'h12: {y00, y01} <= 8'hc9;
    8'h13: {y00, y01} <= 8'h7d;
    8'h14: {y00, y01} <= 8'hfa;
    8'h15: {y00, y01} <= 8'h59;
    8'h16: {y00, y01} <= 8'h47;
    8'h17: {y00, y01} <= 8'hf0;
    8'h18: {y00, y01} <= 8'had;
    8'h19: {y00, y01} <= 8'hd4;
    8'h1a: {y00, y01} <= 8'ha2;
    8'h1b: {y00, y01} <= 8'haf;
    8'h1c: {y00, y01} <= 8'h9c;
    8'h1d: {y00, y01} <= 8'ha4;
    8'h1e: {y00, y01} <= 8'h72;
    8'h1f: {y00, y01} <= 8'hc0;
    8'h20: {y00, y01} <= 8'hb7;
    8'h21: {y00, y01} <= 8'hfd;
    8'h22: {y00, y01} <= 8'h93;
    8'h23: {y00, y01} <= 8'h26;
    8'h24: {y00, y01} <= 8'h36;
    8'h25: {y00, y01} <= 8'h3f;
    8'h26: {y00, y01} <= 8'hf7;
    8'h27: {y00, y01} <= 8'hcc;
    8'h28: {y00, y01} <= 8'h34;
    8'h29: {y00, y01} <= 8'ha5;
    8'h2a: {y00, y01} <= 8'he5;
    8'h2b: {y00, y01} <= 8'hf1;
    8'h2c: {y00, y01} <= 8'h71;
    8'h2d: {y00, y01} <= 8'hd8;
    8'h2e: {y00, y01} <= 8'h31;
    8'h2f: {y00, y01} <= 8'h15;
    8'h30: {y00, y01} <= 8'h04;
    8'h31: {y00, y01} <= 8'hc7;
    8'h32: {y00, y01} <= 8'h23;
    8'h33: {y00, y01} <= 8'hc3;
    8'h34: {y00, y01} <= 8'h18;
    8'h35: {y00, y01} <= 8'h96;
    8'h36: {y00, y01} <= 8'h05;
    8'h37: {y00, y01} <= 8'h9a;
    8'h38: {y00, y01} <= 8'h07;
    8'h39: {y00, y01} <= 8'h12;
    8'h3a: {y00, y01} <= 8'h80;
    8'h3b: {y00, y01} <= 8'he2;
    8'h3c: {y00, y01} <= 8'heb;
    8'h3d: {y00, y01} <= 8'h27;
    8'h3e: {y00, y01} <= 8'hb2;
    8'h3f: {y00, y01} <= 8'h75;
    8'h40: {y00, y01} <= 8'h09;
    8'h41: {y00, y01} <= 8'h83;
    8'h42: {y00, y01} <= 8'h2c;
    8'h43: {y00, y01} <= 8'h1a;
    8'h44: {y00, y01} <= 8'h1b;
    8'h45: {y00, y01} <= 8'h6e;
    8'h46: {y00, y01} <= 8'h5a;
    8'h47: {y00, y01} <= 8'ha0;
    8'h48: {y00, y01} <= 8'h52;
    8'h49: {y00, y01} <= 8'h3b;
    8'h4a: {y00, y01} <= 8'hd6;
    8'h4b: {y00, y01} <= 8'hb3;
    8'h4c: {y00, y01} <= 8'h29;
    8'h4d: {y00, y01} <= 8'he3;
    8'h4e: {y00, y01} <= 8'h2f;
    8'h4f: {y00, y01} <= 8'h84;
    8'h50: {y00, y01} <= 8'h53;
    8'h51: {y00, y01} <= 8'hd1;
    8'h52: {y00, y01} <= 8'h00;
    8'h53: {y00, y01} <= 8'hed;
    8'h54: {y00, y01} <= 8'h20;
    8'h55: {y00, y01} <= 8'hfc;
    8'h56: {y00, y01} <= 8'hb1;
    8'h57: {y00, y01} <= 8'h5b;
    8'h58: {y00, y01} <= 8'h6a;
    8'h59: {y00, y01} <= 8'hcb;
    8'h5a: {y00, y01} <= 8'hbe;
    8'h5b: {y00, y01} <= 8'h39;
    8'h5c: {y00, y01} <= 8'h4a;
    8'h5d: {y00, y01} <= 8'h4c;
    8'h5e: {y00, y01} <= 8'h58;
    8'h5f: {y00, y01} <= 8'hcf;
    8'h60: {y00, y01} <= 8'hd0;
    8'h61: {y00, y01} <= 8'hef;
    8'h62: {y00, y01} <= 8'haa;
    8'h63: {y00, y01} <= 8'hfb;
    8'h64: {y00, y01} <= 8'h43;
    8'h65: {y00, y01} <= 8'h4d;
    8'h66: {y00, y01} <= 8'h33;
    8'h67: {y00, y01} <= 8'h85;
    8'h68: {y00, y01} <= 8'h45;
    8'h69: {y00, y01} <= 8'hf9;
    8'h6a: {y00, y01} <= 8'h02;
    8'h6b: {y00, y01} <= 8'h7f;
    8'h6c: {y00, y01} <= 8'h50;
    8'h6d: {y00, y01} <= 8'h3c;
    8'h6e: {y00, y01} <= 8'h9f;
    8'h6f: {y00, y01} <= 8'ha8;
    8'h70: {y00, y01} <= 8'h51;
    8'h71: {y00, y01} <= 8'ha3;
    8'h72: {y00, y01} <= 8'h40;
    8'h73: {y00, y01} <= 8'h8f;
    8'h74: {y00, y01} <= 8'h92;
    8'h75: {y00, y01} <= 8'h9d;
    8'h76: {y00, y01} <= 8'h38;
    8'h77: {y00, y01} <= 8'hf5;
    8'h78: {y00, y01} <= 8'hbc;
    8'h79: {y00, y01} <= 8'hb6;
    8'h7a: {y00, y01} <= 8'hda;
    8'h7b: {y00, y01} <= 8'h21;
    8'h7c: {y00, y01} <= 8'h10;
    8'h7d: {y00, y01} <= 8'hff;
    8'h7e: {y00, y01} <= 8'hf3;
    8'h7f: {y00, y01} <= 8'hd2;
    8'h80: {y00, y01} <= 8'hcd;
    8'h81: {y00, y01} <= 8'h0c;
    8'h82: {y00, y01} <= 8'h13;
    8'h83: {y00, y01} <= 8'hec;
    8'h84: {y00, y01} <= 8'h5f;
    8'h85: {y00, y01} <= 8'h97;
    8'h86: {y00, y01} <= 8'h44;
    8'h87: {y00, y01} <= 8'h17;
    8'h88: {y00, y01} <= 8'hc4;
    8'h89: {y00, y01} <= 8'ha7;
    8'h8a: {y00, y01} <= 8'h7e;
    8'h8b: {y00, y01} <= 8'h3d;
    8'h8c: {y00, y01} <= 8'h64;
    8'h8d: {y00, y01} <= 8'h5d;
    8'h8e: {y00, y01} <= 8'h19;
    8'h8f: {y00, y01} <= 8'h73;
    8'h90: {y00, y01} <= 8'h60;
    8'h91: {y00, y01} <= 8'h81;
    8'h92: {y00, y01} <= 8'h4f;
    8'h93: {y00, y01} <= 8'hdc;
    8'h94: {y00, y01} <= 8'h22;
    8'h95: {y00, y01} <= 8'h2a;
    8'h96: {y00, y01} <= 8'h90;
    8'h97: {y00, y01} <= 8'h88;
    8'h98: {y00, y01} <= 8'h46;
    8'h99: {y00, y01} <= 8'hee;
    8'h9a: {y00, y01} <= 8'hb8;
    8'h9b: {y00, y01} <= 8'h14;
    8'h9c: {y00, y01} <= 8'hde;
    8'h9d: {y00, y01} <= 8'h5e;
    8'h9e: {y00, y01} <= 8'h0b;
    8'h9f: {y00, y01} <= 8'hdb;
    8'ha0: {y00, y01} <= 8'he0;
    8'ha1: {y00, y01} <= 8'h32;
    8'ha2: {y00, y01} <= 8'h3a;
    8'ha3: {y00, y01} <= 8'h0a;
    8'ha4: {y00, y01} <= 8'h49;
    8'ha5: {y00, y01} <= 8'h06;
    8'ha6: {y00, y01} <= 8'h24;
    8'ha7: {y00, y01} <= 8'h5c;
    8'ha8: {y00, y01} <= 8'hc2;
    8'ha9: {y00, y01} <= 8'hd3;
    8'haa: {y00, y01} <= 8'hac;
    8'hab: {y00, y01} <= 8'h62;
    8'hac: {y00, y01} <= 8'h91;
    8'had: {y00, y01} <= 8'h95;
    8'hae: {y00, y01} <= 8'he4;
    8'haf: {y00, y01} <= 8'h79;
    8'hb0: {y00, y01} <= 8'he7;
    8'hb1: {y00, y01} <= 8'hc8;
    8'hb2: {y00, y01} <= 8'h37;
    8'hb3: {y00, y01} <= 8'h6d;
    8'hb4: {y00, y01} <= 8'h8d;
    8'hb5: {y00, y01} <= 8'hd5;
    8'hb6: {y00, y01} <= 8'h4e;
    8'hb7: {y00, y01} <= 8'ha9;
    8'hb8: {y00, y01} <= 8'h6c;
    8'hb9: {y00, y01} <= 8'h56;
    8'hba: {y00, y01} <= 8'hf4;
    8'hbb: {y00, y01} <= 8'hea;
    8'hbc: {y00, y01} <= 8'h65;
    8'hbd: {y00, y01} <= 8'h7a;
    8'hbe: {y00, y01} <= 8'hae;
    8'hbf: {y00, y01} <= 8'h08;
    8'hc0: {y00, y01} <= 8'hba;
    8'hc1: {y00, y01} <= 8'h78;
    8'hc2: {y00, y01} <= 8'h25;
    8'hc3: {y00, y01} <= 8'h2e;
    8'hc4: {y00, y01} <= 8'h1c;
    8'hc5: {y00, y01} <= 8'ha6;
    8'hc6: {y00, y01} <= 8'hb4;
    8'hc7: {y00, y01} <= 8'hc6;
    8'hc8: {y00, y01} <= 8'he8;
    8'hc9: {y00, y01} <= 8'hdd;
    8'hca: {y00, y01} <= 8'h74;
    8'hcb: {y00, y01} <= 8'h1f;
    8'hcc: {y00, y01} <= 8'h4b;
    8'hcd: {y00, y01} <= 8'hbd;
    8'hce: {y00, y01} <= 8'h8b;
    8'hcf: {y00, y01} <= 8'h8a;
    8'hd0: {y00, y01} <= 8'h70;
    8'hd1: {y00, y01} <= 8'h3e;
    8'hd2: {y00, y01} <= 8'hb5;
    8'hd3: {y00, y01} <= 8'h66;
    8'hd4: {y00, y01} <= 8'h48;
    8'hd5: {y00, y01} <= 8'h03;
    8'hd6: {y00, y01} <= 8'hf6;
    8'hd7: {y00, y01} <= 8'h0e;
    8'hd8: {y00, y01} <= 8'h61;
    8'hd9: {y00, y01} <= 8'h35;
    8'hda: {y00, y01} <= 8'h57;
    8'hdb: {y00, y01} <= 8'hb9;
    8'hdc: {y00, y01} <= 8'h86;
    8'hdd: {y00, y01} <= 8'hc1;
    8'hde: {y00, y01} <= 8'h1d;
    8'hdf: {y00, y01} <= 8'h9e;
    8'he0: {y00, y01} <= 8'he1;
    8'he1: {y00, y01} <= 8'hf8;
    8'he2: {y00, y01} <= 8'h98;
    8'he3: {y00, y01} <= 8'h11;
    8'he4: {y00, y01} <= 8'h69;
    8'he5: {y00, y01} <= 8'hd9;
    8'he6: {y00, y01} <= 8'h8e;
    8'he7: {y00, y01} <= 8'h94;
    8'he8: {y00, y01} <= 8'h9b;
    8'he9: {y00, y01} <= 8'h1e;
    8'hea: {y00, y01} <= 8'h87;
    8'heb: {y00, y01} <= 8'he9;
    8'hec: {y00, y01} <= 8'hce;
    8'hed: {y00, y01} <= 8'h55;
    8'hee: {y00, y01} <= 8'h28;
    8'hef: {y00, y01} <= 8'hdf;
    8'hf0: {y00, y01} <= 8'h8c;
    8'hf1: {y00, y01} <= 8'ha1;
    8'hf2: {y00, y01} <= 8'h89;
    8'hf3: {y00, y01} <= 8'h0d;
    8'hf4: {y00, y01} <= 8'hbf;
    8'hf5: {y00, y01} <= 8'he6;
    8'hf6: {y00, y01} <= 8'h42;
    8'hf7: {y00, y01} <= 8'h68;
    8'hf8: {y00, y01} <= 8'h41;
    8'hf9: {y00, y01} <= 8'h99;
    8'hfa: {y00, y01} <= 8'h2d;
    8'hfb: {y00, y01} <= 8'h0f;
    8'hfc: {y00, y01} <= 8'hb0;
    8'hfd: {y00, y01} <= 8'h54;
    8'hfe: {y00, y01} <= 8'hbb;
    8'hff: {y00, y01} <= 8'h16;
    endcase
	
	
	
	
    // Second Portion
    case (z1)
    8'h00: {y10, y11} <= 8'h63;
    8'h01: {y10, y11} <= 8'h7c;
    8'h02: {y10, y11} <= 8'h77;
    8'h03: {y10, y11} <= 8'h7b;
    8'h04: {y10, y11} <= 8'hf2;
    8'h05: {y10, y11} <= 8'h6b;
    8'h06: {y10, y11} <= 8'h6f;
    8'h07: {y10, y11} <= 8'hc5;
    8'h08: {y10, y11} <= 8'h30;
    8'h09: {y10, y11} <= 8'h01;
    8'h0a: {y10, y11} <= 8'h67;
    8'h0b: {y10, y11} <= 8'h2b;
    8'h0c: {y10, y11} <= 8'hfe;
    8'h0d: {y10, y11} <= 8'hd7;
    8'h0e: {y10, y11} <= 8'hab;
    8'h0f: {y10, y11} <= 8'h76;
    8'h10: {y10, y11} <= 8'hca;
    8'h11: {y10, y11} <= 8'h82;
    8'h12: {y10, y11} <= 8'hc9;
    8'h13: {y10, y11} <= 8'h7d;
    8'h14: {y10, y11} <= 8'hfa;
    8'h15: {y10, y11} <= 8'h59;
    8'h16: {y10, y11} <= 8'h47;
    8'h17: {y10, y11} <= 8'hf0;
    8'h18: {y10, y11} <= 8'had;
    8'h19: {y10, y11} <= 8'hd4;
    8'h1a: {y10, y11} <= 8'ha2;
    8'h1b: {y10, y11} <= 8'haf;
    8'h1c: {y10, y11} <= 8'h9c;
    8'h1d: {y10, y11} <= 8'ha4;
    8'h1e: {y10, y11} <= 8'h72;
    8'h1f: {y10, y11} <= 8'hc0;
    8'h20: {y10, y11} <= 8'hb7;
    8'h21: {y10, y11} <= 8'hfd;
    8'h22: {y10, y11} <= 8'h93;
    8'h23: {y10, y11} <= 8'h26;
    8'h24: {y10, y11} <= 8'h36;
    8'h25: {y10, y11} <= 8'h3f;
    8'h26: {y10, y11} <= 8'hf7;
    8'h27: {y10, y11} <= 8'hcc;
    8'h28: {y10, y11} <= 8'h34;
    8'h29: {y10, y11} <= 8'ha5;
    8'h2a: {y10, y11} <= 8'he5;
    8'h2b: {y10, y11} <= 8'hf1;
    8'h2c: {y10, y11} <= 8'h71;
    8'h2d: {y10, y11} <= 8'hd8;
    8'h2e: {y10, y11} <= 8'h31;
    8'h2f: {y10, y11} <= 8'h15;
    8'h30: {y10, y11} <= 8'h04;
    8'h31: {y10, y11} <= 8'hc7;
    8'h32: {y10, y11} <= 8'h23;
    8'h33: {y10, y11} <= 8'hc3;
    8'h34: {y10, y11} <= 8'h18;
    8'h35: {y10, y11} <= 8'h96;
    8'h36: {y10, y11} <= 8'h05;
    8'h37: {y10, y11} <= 8'h9a;
    8'h38: {y10, y11} <= 8'h07;
    8'h39: {y10, y11} <= 8'h12;
    8'h3a: {y10, y11} <= 8'h80;
    8'h3b: {y10, y11} <= 8'he2;
    8'h3c: {y10, y11} <= 8'heb;
    8'h3d: {y10, y11} <= 8'h27;
    8'h3e: {y10, y11} <= 8'hb2;
    8'h3f: {y10, y11} <= 8'h75;
    8'h40: {y10, y11} <= 8'h09;
    8'h41: {y10, y11} <= 8'h83;
    8'h42: {y10, y11} <= 8'h2c;
    8'h43: {y10, y11} <= 8'h1a;
    8'h44: {y10, y11} <= 8'h1b;
    8'h45: {y10, y11} <= 8'h6e;
    8'h46: {y10, y11} <= 8'h5a;
    8'h47: {y10, y11} <= 8'ha0;
    8'h48: {y10, y11} <= 8'h52;
    8'h49: {y10, y11} <= 8'h3b;
    8'h4a: {y10, y11} <= 8'hd6;
    8'h4b: {y10, y11} <= 8'hb3;
    8'h4c: {y10, y11} <= 8'h29;
    8'h4d: {y10, y11} <= 8'he3;
    8'h4e: {y10, y11} <= 8'h2f;
    8'h4f: {y10, y11} <= 8'h84;
    8'h50: {y10, y11} <= 8'h53;
    8'h51: {y10, y11} <= 8'hd1;
    8'h52: {y10, y11} <= 8'h00;
    8'h53: {y10, y11} <= 8'hed;
    8'h54: {y10, y11} <= 8'h20;
    8'h55: {y10, y11} <= 8'hfc;
    8'h56: {y10, y11} <= 8'hb1;
    8'h57: {y10, y11} <= 8'h5b;
    8'h58: {y10, y11} <= 8'h6a;
    8'h59: {y10, y11} <= 8'hcb;
    8'h5a: {y10, y11} <= 8'hbe;
    8'h5b: {y10, y11} <= 8'h39;
    8'h5c: {y10, y11} <= 8'h4a;
    8'h5d: {y10, y11} <= 8'h4c;
    8'h5e: {y10, y11} <= 8'h58;
    8'h5f: {y10, y11} <= 8'hcf;
    8'h60: {y10, y11} <= 8'hd0;
    8'h61: {y10, y11} <= 8'hef;
    8'h62: {y10, y11} <= 8'haa;
    8'h63: {y10, y11} <= 8'hfb;
    8'h64: {y10, y11} <= 8'h43;
    8'h65: {y10, y11} <= 8'h4d;
    8'h66: {y10, y11} <= 8'h33;
    8'h67: {y10, y11} <= 8'h85;
    8'h68: {y10, y11} <= 8'h45;
    8'h69: {y10, y11} <= 8'hf9;
    8'h6a: {y10, y11} <= 8'h02;
    8'h6b: {y10, y11} <= 8'h7f;
    8'h6c: {y10, y11} <= 8'h50;
    8'h6d: {y10, y11} <= 8'h3c;
    8'h6e: {y10, y11} <= 8'h9f;
    8'h6f: {y10, y11} <= 8'ha8;
    8'h70: {y10, y11} <= 8'h51;
    8'h71: {y10, y11} <= 8'ha3;
    8'h72: {y10, y11} <= 8'h40;
    8'h73: {y10, y11} <= 8'h8f;
    8'h74: {y10, y11} <= 8'h92;
    8'h75: {y10, y11} <= 8'h9d;
    8'h76: {y10, y11} <= 8'h38;
    8'h77: {y10, y11} <= 8'hf5;
    8'h78: {y10, y11} <= 8'hbc;
    8'h79: {y10, y11} <= 8'hb6;
    8'h7a: {y10, y11} <= 8'hda;
    8'h7b: {y10, y11} <= 8'h21;
    8'h7c: {y10, y11} <= 8'h10;
    8'h7d: {y10, y11} <= 8'hff;
    8'h7e: {y10, y11} <= 8'hf3;
    8'h7f: {y10, y11} <= 8'hd2;
    8'h80: {y10, y11} <= 8'hcd;
    8'h81: {y10, y11} <= 8'h0c;
    8'h82: {y10, y11} <= 8'h13;
    8'h83: {y10, y11} <= 8'hec;
    8'h84: {y10, y11} <= 8'h5f;
    8'h85: {y10, y11} <= 8'h97;
    8'h86: {y10, y11} <= 8'h44;
    8'h87: {y10, y11} <= 8'h17;
    8'h88: {y10, y11} <= 8'hc4;
    8'h89: {y10, y11} <= 8'ha7;
    8'h8a: {y10, y11} <= 8'h7e;
    8'h8b: {y10, y11} <= 8'h3d;
    8'h8c: {y10, y11} <= 8'h64;
    8'h8d: {y10, y11} <= 8'h5d;
    8'h8e: {y10, y11} <= 8'h19;
    8'h8f: {y10, y11} <= 8'h73;
    8'h90: {y10, y11} <= 8'h60;
    8'h91: {y10, y11} <= 8'h81;
    8'h92: {y10, y11} <= 8'h4f;
    8'h93: {y10, y11} <= 8'hdc;
    8'h94: {y10, y11} <= 8'h22;
    8'h95: {y10, y11} <= 8'h2a;
    8'h96: {y10, y11} <= 8'h90;
    8'h97: {y10, y11} <= 8'h88;
    8'h98: {y10, y11} <= 8'h46;
    8'h99: {y10, y11} <= 8'hee;
    8'h9a: {y10, y11} <= 8'hb8;
    8'h9b: {y10, y11} <= 8'h14;
    8'h9c: {y10, y11} <= 8'hde;
    8'h9d: {y10, y11} <= 8'h5e;
    8'h9e: {y10, y11} <= 8'h0b;
    8'h9f: {y10, y11} <= 8'hdb;
    8'ha0: {y10, y11} <= 8'he0;
    8'ha1: {y10, y11} <= 8'h32;
    8'ha2: {y10, y11} <= 8'h3a;
    8'ha3: {y10, y11} <= 8'h0a;
    8'ha4: {y10, y11} <= 8'h49;
    8'ha5: {y10, y11} <= 8'h06;
    8'ha6: {y10, y11} <= 8'h24;
    8'ha7: {y10, y11} <= 8'h5c;
    8'ha8: {y10, y11} <= 8'hc2;
    8'ha9: {y10, y11} <= 8'hd3;
    8'haa: {y10, y11} <= 8'hac;
    8'hab: {y10, y11} <= 8'h62;
    8'hac: {y10, y11} <= 8'h91;
    8'had: {y10, y11} <= 8'h95;
    8'hae: {y10, y11} <= 8'he4;
    8'haf: {y10, y11} <= 8'h79;
    8'hb0: {y10, y11} <= 8'he7;
    8'hb1: {y10, y11} <= 8'hc8;
    8'hb2: {y10, y11} <= 8'h37;
    8'hb3: {y10, y11} <= 8'h6d;
    8'hb4: {y10, y11} <= 8'h8d;
    8'hb5: {y10, y11} <= 8'hd5;
    8'hb6: {y10, y11} <= 8'h4e;
    8'hb7: {y10, y11} <= 8'ha9;
    8'hb8: {y10, y11} <= 8'h6c;
    8'hb9: {y10, y11} <= 8'h56;
    8'hba: {y10, y11} <= 8'hf4;
    8'hbb: {y10, y11} <= 8'hea;
    8'hbc: {y10, y11} <= 8'h65;
    8'hbd: {y10, y11} <= 8'h7a;
    8'hbe: {y10, y11} <= 8'hae;
    8'hbf: {y10, y11} <= 8'h08;
    8'hc0: {y10, y11} <= 8'hba;
    8'hc1: {y10, y11} <= 8'h78;
    8'hc2: {y10, y11} <= 8'h25;
    8'hc3: {y10, y11} <= 8'h2e;
    8'hc4: {y10, y11} <= 8'h1c;
    8'hc5: {y10, y11} <= 8'ha6;
    8'hc6: {y10, y11} <= 8'hb4;
    8'hc7: {y10, y11} <= 8'hc6;
    8'hc8: {y10, y11} <= 8'he8;
    8'hc9: {y10, y11} <= 8'hdd;
    8'hca: {y10, y11} <= 8'h74;
    8'hcb: {y10, y11} <= 8'h1f;
    8'hcc: {y10, y11} <= 8'h4b;
    8'hcd: {y10, y11} <= 8'hbd;
    8'hce: {y10, y11} <= 8'h8b;
    8'hcf: {y10, y11} <= 8'h8a;
    8'hd0: {y10, y11} <= 8'h70;
    8'hd1: {y10, y11} <= 8'h3e;
    8'hd2: {y10, y11} <= 8'hb5;
    8'hd3: {y10, y11} <= 8'h66;
    8'hd4: {y10, y11} <= 8'h48;
    8'hd5: {y10, y11} <= 8'h03;
    8'hd6: {y10, y11} <= 8'hf6;
    8'hd7: {y10, y11} <= 8'h0e;
    8'hd8: {y10, y11} <= 8'h61;
    8'hd9: {y10, y11} <= 8'h35;
    8'hda: {y10, y11} <= 8'h57;
    8'hdb: {y10, y11} <= 8'hb9;
    8'hdc: {y10, y11} <= 8'h86;
    8'hdd: {y10, y11} <= 8'hc1;
    8'hde: {y10, y11} <= 8'h1d;
    8'hdf: {y10, y11} <= 8'h9e;
    8'he0: {y10, y11} <= 8'he1;
    8'he1: {y10, y11} <= 8'hf8;
    8'he2: {y10, y11} <= 8'h98;
    8'he3: {y10, y11} <= 8'h11;
    8'he4: {y10, y11} <= 8'h69;
    8'he5: {y10, y11} <= 8'hd9;
    8'he6: {y10, y11} <= 8'h8e;
    8'he7: {y10, y11} <= 8'h94;
    8'he8: {y10, y11} <= 8'h9b;
    8'he9: {y10, y11} <= 8'h1e;
    8'hea: {y10, y11} <= 8'h87;
    8'heb: {y10, y11} <= 8'he9;
    8'hec: {y10, y11} <= 8'hce;
    8'hed: {y10, y11} <= 8'h55;
    8'hee: {y10, y11} <= 8'h28;
    8'hef: {y10, y11} <= 8'hdf;
    8'hf0: {y10, y11} <= 8'h8c;
    8'hf1: {y10, y11} <= 8'ha1;
    8'hf2: {y10, y11} <= 8'h89;
    8'hf3: {y10, y11} <= 8'h0d;
    8'hf4: {y10, y11} <= 8'hbf;
    8'hf5: {y10, y11} <= 8'he6;
    8'hf6: {y10, y11} <= 8'h42;
    8'hf7: {y10, y11} <= 8'h68;
    8'hf8: {y10, y11} <= 8'h41;
    8'hf9: {y10, y11} <= 8'h99;
    8'hfa: {y10, y11} <= 8'h2d;
    8'hfb: {y10, y11} <= 8'h0f;
    8'hfc: {y10, y11} <= 8'hb0;
    8'hfd: {y10, y11} <= 8'h54;
    8'hfe: {y10, y11} <= 8'hbb;
    8'hff: {y10, y11} <= 8'h16;
    endcase
	
    end
	
    assign g0 = {y00, y11} ^ k0_o;
    assign g1 = {y10, y01} ^ k1_o;

    always @ (posedge clk) begin
        out <= {g0, g1};
    end

endmodule
